// Benchmark "C1355.iscas" written by ABC on Thu Mar 19 13:02:35 2020

module C1355_iscas  ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31;
  wire new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_,
    new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_,
    new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_,
    new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_, new_n111_, new_n112_, new_n113_,
    new_n114_, new_n115_, new_n116_, new_n117_, new_n118_, new_n119_,
    new_n120_, new_n121_, new_n122_, new_n123_, new_n124_, new_n125_,
    new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_,
    new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_;
  assign new_n74_ = pi39 & pi40;
  assign new_n75_ = pi38 & pi40;
  assign new_n76_ = pi37 & pi40;
  assign new_n77_ = pi36 & pi40;
  assign new_n78_ = pi35 & pi40;
  assign new_n79_ = pi34 & pi40;
  assign new_n80_ = pi33 & pi40;
  assign new_n81_ = pi32 & pi40;
  assign new_n82_ = ~pi30 | ~pi31;
  assign new_n83_ = ~pi28 | ~pi29;
  assign new_n84_ = ~pi27 | ~pi31;
  assign new_n85_ = ~pi26 | ~pi30;
  assign new_n86_ = ~pi26 | ~pi27;
  assign new_n87_ = ~pi25 | ~pi29;
  assign new_n88_ = ~pi24 | ~pi28;
  assign new_n89_ = ~pi24 | ~pi25;
  assign new_n90_ = ~pi22 | ~pi23;
  assign new_n91_ = ~pi20 | ~pi21;
  assign new_n92_ = ~pi19 | ~pi23;
  assign new_n93_ = ~pi18 | ~pi22;
  assign new_n94_ = ~pi18 | ~pi19;
  assign new_n95_ = ~pi17 | ~pi21;
  assign new_n96_ = ~pi16 | ~pi20;
  assign new_n97_ = ~pi16 | ~pi17;
  assign new_n98_ = ~pi14 | ~pi15;
  assign new_n99_ = ~pi12 | ~pi13;
  assign new_n100_ = ~pi11 | ~pi15;
  assign new_n101_ = ~pi10 | ~pi14;
  assign new_n102_ = ~pi10 | ~pi11;
  assign new_n103_ = ~pi09 | ~pi13;
  assign new_n104_ = ~pi08 | ~pi12;
  assign new_n105_ = ~pi08 | ~pi09;
  assign new_n106_ = ~pi06 | ~pi07;
  assign new_n107_ = ~pi04 | ~pi05;
  assign new_n108_ = ~pi03 | ~pi07;
  assign new_n109_ = ~pi02 | ~pi06;
  assign new_n110_ = ~pi02 | ~pi03;
  assign new_n111_ = ~pi01 | ~pi05;
  assign new_n112_ = ~pi00 | ~pi04;
  assign new_n113_ = ~pi00 | ~pi01;
  assign new_n114_ = ~pi31 | ~new_n84_;
  assign new_n115_ = ~pi31 | ~new_n82_;
  assign new_n116_ = ~pi30 | ~new_n85_;
  assign new_n117_ = ~pi30 | ~new_n82_;
  assign new_n118_ = ~pi29 | ~new_n87_;
  assign new_n119_ = ~pi29 | ~new_n83_;
  assign new_n120_ = ~pi28 | ~new_n88_;
  assign new_n121_ = ~pi28 | ~new_n83_;
  assign new_n122_ = ~pi27 | ~new_n84_;
  assign new_n123_ = ~pi27 | ~new_n86_;
  assign new_n124_ = ~pi26 | ~new_n85_;
  assign new_n125_ = ~pi26 | ~new_n86_;
  assign new_n126_ = ~pi25 | ~new_n87_;
  assign new_n127_ = ~pi25 | ~new_n89_;
  assign new_n128_ = ~pi24 | ~new_n88_;
  assign new_n129_ = ~pi24 | ~new_n89_;
  assign new_n130_ = ~pi23 | ~new_n92_;
  assign new_n131_ = ~pi23 | ~new_n90_;
  assign new_n132_ = ~pi22 | ~new_n93_;
  assign new_n133_ = ~pi22 | ~new_n90_;
  assign new_n134_ = ~pi21 | ~new_n95_;
  assign new_n135_ = ~pi21 | ~new_n91_;
  assign new_n136_ = ~pi20 | ~new_n96_;
  assign new_n137_ = ~pi20 | ~new_n91_;
  assign new_n138_ = ~pi19 | ~new_n92_;
  assign new_n139_ = ~pi19 | ~new_n94_;
  assign new_n140_ = ~pi18 | ~new_n93_;
  assign new_n141_ = ~pi18 | ~new_n94_;
  assign new_n142_ = ~pi17 | ~new_n95_;
  assign new_n143_ = ~pi17 | ~new_n97_;
  assign new_n144_ = ~pi16 | ~new_n96_;
  assign new_n145_ = ~pi16 | ~new_n97_;
  assign new_n146_ = ~pi15 | ~new_n100_;
  assign new_n147_ = ~pi15 | ~new_n98_;
  assign new_n148_ = ~pi14 | ~new_n101_;
  assign new_n149_ = ~pi14 | ~new_n98_;
  assign new_n150_ = ~pi13 | ~new_n103_;
  assign new_n151_ = ~pi13 | ~new_n99_;
  assign new_n152_ = ~pi12 | ~new_n104_;
  assign new_n153_ = ~pi12 | ~new_n99_;
  assign new_n154_ = ~pi11 | ~new_n100_;
  assign new_n155_ = ~pi11 | ~new_n102_;
  assign new_n156_ = ~pi10 | ~new_n101_;
  assign new_n157_ = ~pi10 | ~new_n102_;
  assign new_n158_ = ~pi09 | ~new_n103_;
  assign new_n159_ = ~pi09 | ~new_n105_;
  assign new_n160_ = ~pi08 | ~new_n104_;
  assign new_n161_ = ~pi08 | ~new_n105_;
  assign new_n162_ = ~pi07 | ~new_n108_;
  assign new_n163_ = ~pi07 | ~new_n106_;
  assign new_n164_ = ~pi06 | ~new_n109_;
  assign new_n165_ = ~pi06 | ~new_n106_;
  assign new_n166_ = ~pi05 | ~new_n111_;
  assign new_n167_ = ~pi05 | ~new_n107_;
  assign new_n168_ = ~pi04 | ~new_n112_;
  assign new_n169_ = ~pi04 | ~new_n107_;
  assign new_n170_ = ~pi03 | ~new_n108_;
  assign new_n171_ = ~pi03 | ~new_n110_;
  assign new_n172_ = ~pi02 | ~new_n109_;
  assign new_n173_ = ~pi02 | ~new_n110_;
  assign new_n174_ = ~pi01 | ~new_n111_;
  assign new_n175_ = ~pi01 | ~new_n113_;
  assign new_n176_ = ~pi00 | ~new_n112_;
  assign new_n177_ = ~pi00 | ~new_n113_;
  assign new_n178_ = ~new_n122_ | ~new_n114_;
  assign new_n179_ = ~new_n117_ | ~new_n115_;
  assign new_n180_ = ~new_n124_ | ~new_n116_;
  assign new_n181_ = ~new_n126_ | ~new_n118_;
  assign new_n182_ = ~new_n121_ | ~new_n119_;
  assign new_n183_ = ~new_n128_ | ~new_n120_;
  assign new_n184_ = ~new_n125_ | ~new_n123_;
  assign new_n185_ = ~new_n129_ | ~new_n127_;
  assign new_n186_ = ~new_n138_ | ~new_n130_;
  assign new_n187_ = ~new_n133_ | ~new_n131_;
  assign new_n188_ = ~new_n140_ | ~new_n132_;
  assign new_n189_ = ~new_n142_ | ~new_n134_;
  assign new_n190_ = ~new_n137_ | ~new_n135_;
  assign new_n191_ = ~new_n144_ | ~new_n136_;
  assign new_n192_ = ~new_n141_ | ~new_n139_;
  assign new_n193_ = ~new_n145_ | ~new_n143_;
  assign new_n194_ = ~new_n154_ | ~new_n146_;
  assign new_n195_ = ~new_n149_ | ~new_n147_;
  assign new_n196_ = ~new_n156_ | ~new_n148_;
  assign new_n197_ = ~new_n158_ | ~new_n150_;
  assign new_n198_ = ~new_n153_ | ~new_n151_;
  assign new_n199_ = ~new_n160_ | ~new_n152_;
  assign new_n200_ = ~new_n157_ | ~new_n155_;
  assign new_n201_ = ~new_n161_ | ~new_n159_;
  assign new_n202_ = ~new_n170_ | ~new_n162_;
  assign new_n203_ = ~new_n165_ | ~new_n163_;
  assign new_n204_ = ~new_n172_ | ~new_n164_;
  assign new_n205_ = ~new_n174_ | ~new_n166_;
  assign new_n206_ = ~new_n169_ | ~new_n167_;
  assign new_n207_ = ~new_n176_ | ~new_n168_;
  assign new_n208_ = ~new_n173_ | ~new_n171_;
  assign new_n209_ = ~new_n177_ | ~new_n175_;
  assign new_n210_ = ~new_n186_ | ~new_n178_;
  assign new_n211_ = ~new_n182_ | ~new_n179_;
  assign new_n212_ = ~new_n188_ | ~new_n180_;
  assign new_n213_ = ~new_n189_ | ~new_n181_;
  assign new_n214_ = ~new_n191_ | ~new_n183_;
  assign new_n215_ = ~new_n185_ | ~new_n184_;
  assign new_n216_ = ~new_n190_ | ~new_n187_;
  assign new_n217_ = ~new_n193_ | ~new_n192_;
  assign new_n218_ = ~new_n202_ | ~new_n194_;
  assign new_n219_ = ~new_n198_ | ~new_n195_;
  assign new_n220_ = ~new_n204_ | ~new_n196_;
  assign new_n221_ = ~new_n205_ | ~new_n197_;
  assign new_n222_ = ~new_n207_ | ~new_n199_;
  assign new_n223_ = ~new_n201_ | ~new_n200_;
  assign new_n224_ = ~new_n206_ | ~new_n203_;
  assign new_n225_ = ~new_n209_ | ~new_n208_;
  assign new_n226_ = ~new_n178_ | ~new_n210_;
  assign new_n227_ = ~new_n179_ | ~new_n211_;
  assign new_n228_ = ~new_n180_ | ~new_n212_;
  assign new_n229_ = ~new_n181_ | ~new_n213_;
  assign new_n230_ = ~new_n182_ | ~new_n211_;
  assign new_n231_ = ~new_n183_ | ~new_n214_;
  assign new_n232_ = ~new_n184_ | ~new_n215_;
  assign new_n233_ = ~new_n185_ | ~new_n215_;
  assign new_n234_ = ~new_n186_ | ~new_n210_;
  assign new_n235_ = ~new_n187_ | ~new_n216_;
  assign new_n236_ = ~new_n188_ | ~new_n212_;
  assign new_n237_ = ~new_n189_ | ~new_n213_;
  assign new_n238_ = ~new_n190_ | ~new_n216_;
  assign new_n239_ = ~new_n191_ | ~new_n214_;
  assign new_n240_ = ~new_n192_ | ~new_n217_;
  assign new_n241_ = ~new_n193_ | ~new_n217_;
  assign new_n242_ = ~new_n194_ | ~new_n218_;
  assign new_n243_ = ~new_n195_ | ~new_n219_;
  assign new_n244_ = ~new_n196_ | ~new_n220_;
  assign new_n245_ = ~new_n197_ | ~new_n221_;
  assign new_n246_ = ~new_n198_ | ~new_n219_;
  assign new_n247_ = ~new_n199_ | ~new_n222_;
  assign new_n248_ = ~new_n200_ | ~new_n223_;
  assign new_n249_ = ~new_n201_ | ~new_n223_;
  assign new_n250_ = ~new_n202_ | ~new_n218_;
  assign new_n251_ = ~new_n203_ | ~new_n224_;
  assign new_n252_ = ~new_n204_ | ~new_n220_;
  assign new_n253_ = ~new_n205_ | ~new_n221_;
  assign new_n254_ = ~new_n206_ | ~new_n224_;
  assign new_n255_ = ~new_n207_ | ~new_n222_;
  assign new_n256_ = ~new_n208_ | ~new_n225_;
  assign new_n257_ = ~new_n209_ | ~new_n225_;
  assign new_n258_ = ~new_n234_ | ~new_n226_;
  assign new_n259_ = ~new_n230_ | ~new_n227_;
  assign new_n260_ = ~new_n236_ | ~new_n228_;
  assign new_n261_ = ~new_n237_ | ~new_n229_;
  assign new_n262_ = ~new_n239_ | ~new_n231_;
  assign new_n263_ = ~new_n233_ | ~new_n232_;
  assign new_n264_ = ~new_n238_ | ~new_n235_;
  assign new_n265_ = ~new_n241_ | ~new_n240_;
  assign new_n266_ = ~new_n250_ | ~new_n242_;
  assign new_n267_ = ~new_n246_ | ~new_n243_;
  assign new_n268_ = ~new_n252_ | ~new_n244_;
  assign new_n269_ = ~new_n253_ | ~new_n245_;
  assign new_n270_ = ~new_n255_ | ~new_n247_;
  assign new_n271_ = ~new_n249_ | ~new_n248_;
  assign new_n272_ = ~new_n254_ | ~new_n251_;
  assign new_n273_ = ~new_n257_ | ~new_n256_;
  assign new_n274_ = ~new_n263_ | ~new_n259_;
  assign new_n275_ = ~new_n264_ | ~new_n259_;
  assign new_n276_ = ~new_n265_ | ~new_n263_;
  assign new_n277_ = ~new_n265_ | ~new_n264_;
  assign new_n278_ = ~new_n271_ | ~new_n267_;
  assign new_n279_ = ~new_n272_ | ~new_n267_;
  assign new_n280_ = ~new_n273_ | ~new_n271_;
  assign new_n281_ = ~new_n273_ | ~new_n272_;
  assign new_n282_ = ~new_n259_ | ~new_n274_;
  assign new_n283_ = ~new_n259_ | ~new_n275_;
  assign new_n284_ = ~new_n263_ | ~new_n274_;
  assign new_n285_ = ~new_n263_ | ~new_n276_;
  assign new_n286_ = ~new_n264_ | ~new_n277_;
  assign new_n287_ = ~new_n264_ | ~new_n275_;
  assign new_n288_ = ~new_n265_ | ~new_n277_;
  assign new_n289_ = ~new_n265_ | ~new_n276_;
  assign new_n290_ = ~new_n267_ | ~new_n278_;
  assign new_n291_ = ~new_n267_ | ~new_n279_;
  assign new_n292_ = ~new_n271_ | ~new_n278_;
  assign new_n293_ = ~new_n271_ | ~new_n280_;
  assign new_n294_ = ~new_n272_ | ~new_n281_;
  assign new_n295_ = ~new_n272_ | ~new_n279_;
  assign new_n296_ = ~new_n273_ | ~new_n281_;
  assign new_n297_ = ~new_n273_ | ~new_n280_;
  assign new_n298_ = ~new_n284_ | ~new_n282_;
  assign new_n299_ = ~new_n287_ | ~new_n283_;
  assign new_n300_ = ~new_n289_ | ~new_n285_;
  assign new_n301_ = ~new_n288_ | ~new_n286_;
  assign new_n302_ = ~new_n292_ | ~new_n290_;
  assign new_n303_ = ~new_n295_ | ~new_n291_;
  assign new_n304_ = ~new_n297_ | ~new_n293_;
  assign new_n305_ = ~new_n296_ | ~new_n294_;
  assign new_n306_ = ~new_n74_ | ~new_n303_;
  assign new_n307_ = ~new_n75_ | ~new_n304_;
  assign new_n308_ = ~new_n76_ | ~new_n302_;
  assign new_n309_ = ~new_n77_ | ~new_n305_;
  assign new_n310_ = ~new_n78_ | ~new_n299_;
  assign new_n311_ = ~new_n79_ | ~new_n300_;
  assign new_n312_ = ~new_n80_ | ~new_n298_;
  assign new_n313_ = ~new_n81_ | ~new_n301_;
  assign new_n314_ = ~new_n74_ | ~new_n306_;
  assign new_n315_ = ~new_n75_ | ~new_n307_;
  assign new_n316_ = ~new_n76_ | ~new_n308_;
  assign new_n317_ = ~new_n77_ | ~new_n309_;
  assign new_n318_ = ~new_n78_ | ~new_n310_;
  assign new_n319_ = ~new_n79_ | ~new_n311_;
  assign new_n320_ = ~new_n80_ | ~new_n312_;
  assign new_n321_ = ~new_n81_ | ~new_n313_;
  assign new_n322_ = ~new_n298_ | ~new_n312_;
  assign new_n323_ = ~new_n299_ | ~new_n310_;
  assign new_n324_ = ~new_n300_ | ~new_n311_;
  assign new_n325_ = ~new_n301_ | ~new_n313_;
  assign new_n326_ = ~new_n302_ | ~new_n308_;
  assign new_n327_ = ~new_n303_ | ~new_n306_;
  assign new_n328_ = ~new_n304_ | ~new_n307_;
  assign new_n329_ = ~new_n305_ | ~new_n309_;
  assign new_n330_ = ~new_n314_ | ~new_n327_;
  assign new_n331_ = ~new_n315_ | ~new_n328_;
  assign new_n332_ = ~new_n316_ | ~new_n326_;
  assign new_n333_ = ~new_n317_ | ~new_n329_;
  assign new_n334_ = ~new_n318_ | ~new_n323_;
  assign new_n335_ = ~new_n319_ | ~new_n324_;
  assign new_n336_ = ~new_n320_ | ~new_n322_;
  assign new_n337_ = ~new_n321_ | ~new_n325_;
  assign new_n338_ = ~new_n258_ | ~new_n330_;
  assign new_n339_ = ~new_n260_ | ~new_n331_;
  assign new_n340_ = ~new_n261_ | ~new_n332_;
  assign new_n341_ = ~new_n262_ | ~new_n333_;
  assign new_n342_ = ~new_n266_ | ~new_n334_;
  assign new_n343_ = ~new_n268_ | ~new_n335_;
  assign new_n344_ = ~new_n269_ | ~new_n336_;
  assign new_n345_ = ~new_n270_ | ~new_n337_;
  assign new_n346_ = ~new_n330_ | ~new_n338_;
  assign new_n347_ = ~new_n331_ | ~new_n339_;
  assign new_n348_ = ~new_n332_ | ~new_n340_;
  assign new_n349_ = ~new_n333_ | ~new_n341_;
  assign new_n350_ = ~new_n334_ | ~new_n342_;
  assign new_n351_ = ~new_n335_ | ~new_n343_;
  assign new_n352_ = ~new_n336_ | ~new_n344_;
  assign new_n353_ = ~new_n337_ | ~new_n345_;
  assign new_n354_ = ~new_n258_ | ~new_n338_;
  assign new_n355_ = ~new_n260_ | ~new_n339_;
  assign new_n356_ = ~new_n261_ | ~new_n340_;
  assign new_n357_ = ~new_n262_ | ~new_n341_;
  assign new_n358_ = ~new_n266_ | ~new_n342_;
  assign new_n359_ = ~new_n268_ | ~new_n343_;
  assign new_n360_ = ~new_n269_ | ~new_n344_;
  assign new_n361_ = ~new_n270_ | ~new_n345_;
  assign new_n362_ = ~new_n354_ | ~new_n346_;
  assign new_n363_ = ~new_n355_ | ~new_n347_;
  assign new_n364_ = ~new_n356_ | ~new_n348_;
  assign new_n365_ = ~new_n357_ | ~new_n349_;
  assign new_n366_ = ~new_n358_ | ~new_n350_;
  assign new_n367_ = ~new_n359_ | ~new_n351_;
  assign new_n368_ = ~new_n360_ | ~new_n352_;
  assign new_n369_ = ~new_n361_ | ~new_n353_;
  assign new_n370_ = ~new_n362_;
  assign new_n371_ = ~new_n362_;
  assign new_n372_ = ~new_n362_;
  assign new_n373_ = ~new_n362_;
  assign new_n374_ = ~new_n362_;
  assign new_n375_ = ~new_n363_;
  assign new_n376_ = ~new_n363_;
  assign new_n377_ = ~new_n363_;
  assign new_n378_ = ~new_n363_;
  assign new_n379_ = ~new_n363_;
  assign new_n380_ = ~new_n364_;
  assign new_n381_ = ~new_n364_;
  assign new_n382_ = ~new_n364_;
  assign new_n383_ = ~new_n364_;
  assign new_n384_ = ~new_n364_;
  assign new_n385_ = ~new_n365_;
  assign new_n386_ = ~new_n365_;
  assign new_n387_ = ~new_n365_;
  assign new_n388_ = ~new_n365_;
  assign new_n389_ = ~new_n365_;
  assign new_n390_ = ~new_n366_;
  assign new_n391_ = ~new_n366_;
  assign new_n392_ = ~new_n366_;
  assign new_n393_ = ~new_n366_;
  assign new_n394_ = ~new_n366_;
  assign new_n395_ = ~new_n367_;
  assign new_n396_ = ~new_n367_;
  assign new_n397_ = ~new_n367_;
  assign new_n398_ = ~new_n367_;
  assign new_n399_ = ~new_n367_;
  assign new_n400_ = ~new_n368_;
  assign new_n401_ = ~new_n368_;
  assign new_n402_ = ~new_n368_;
  assign new_n403_ = ~new_n368_;
  assign new_n404_ = ~new_n368_;
  assign new_n405_ = ~new_n369_;
  assign new_n406_ = ~new_n369_;
  assign new_n407_ = ~new_n369_;
  assign new_n408_ = ~new_n369_;
  assign new_n409_ = ~new_n369_;
  assign new_n410_ = new_n362_ & new_n377_ & new_n387_ & new_n382_;
  assign new_n411_ = new_n372_ & new_n363_ & new_n388_ & new_n383_;
  assign new_n412_ = new_n373_ & new_n378_ & new_n389_ & new_n364_;
  assign new_n413_ = new_n374_ & new_n379_ & new_n365_ & new_n384_;
  assign new_n414_ = new_n366_ & new_n395_ & new_n405_ & new_n400_;
  assign new_n415_ = new_n390_ & new_n367_ & new_n406_ & new_n401_;
  assign new_n416_ = new_n391_ & new_n396_ & new_n407_ & new_n368_;
  assign new_n417_ = new_n392_ & new_n397_ & new_n369_ & new_n402_;
  assign new_n418_ = new_n413_ | new_n412_ | new_n410_ | new_n411_;
  assign new_n419_ = new_n417_ | new_n416_ | new_n414_ | new_n415_;
  assign new_n420_ = new_n419_ & new_n362_ & new_n375_ & new_n365_ & new_n381_;
  assign new_n421_ = new_n419_ & new_n362_ & new_n376_ & new_n386_ & new_n364_;
  assign new_n422_ = new_n419_ & new_n370_ & new_n363_ & new_n365_ & new_n380_;
  assign new_n423_ = new_n419_ & new_n371_ & new_n363_ & new_n385_ & new_n364_;
  assign new_n424_ = new_n418_ & new_n366_ & new_n398_ & new_n369_ & new_n404_;
  assign new_n425_ = new_n418_ & new_n366_ & new_n399_ & new_n409_ & new_n368_;
  assign new_n426_ = new_n418_ & new_n393_ & new_n367_ & new_n369_ & new_n403_;
  assign new_n427_ = new_n418_ & new_n394_ & new_n367_ & new_n408_ & new_n368_;
  assign new_n428_ = new_n362_ & new_n426_;
  assign new_n429_ = new_n362_ & new_n424_;
  assign new_n430_ = new_n362_ & new_n427_;
  assign new_n431_ = new_n362_ & new_n425_;
  assign new_n432_ = new_n363_ & new_n426_;
  assign new_n433_ = new_n363_ & new_n424_;
  assign new_n434_ = new_n363_ & new_n427_;
  assign new_n435_ = new_n363_ & new_n425_;
  assign new_n436_ = new_n364_ & new_n426_;
  assign new_n437_ = new_n364_ & new_n424_;
  assign new_n438_ = new_n364_ & new_n427_;
  assign new_n439_ = new_n364_ & new_n425_;
  assign new_n440_ = new_n365_ & new_n426_;
  assign new_n441_ = new_n365_ & new_n424_;
  assign new_n442_ = new_n365_ & new_n427_;
  assign new_n443_ = new_n365_ & new_n425_;
  assign new_n444_ = new_n366_ & new_n422_;
  assign new_n445_ = new_n366_ & new_n420_;
  assign new_n446_ = new_n366_ & new_n423_;
  assign new_n447_ = new_n366_ & new_n421_;
  assign new_n448_ = new_n367_ & new_n422_;
  assign new_n449_ = new_n367_ & new_n420_;
  assign new_n450_ = new_n367_ & new_n423_;
  assign new_n451_ = new_n367_ & new_n421_;
  assign new_n452_ = new_n368_ & new_n422_;
  assign new_n453_ = new_n368_ & new_n420_;
  assign new_n454_ = new_n368_ & new_n423_;
  assign new_n455_ = new_n368_ & new_n421_;
  assign new_n456_ = new_n369_ & new_n422_;
  assign new_n457_ = new_n369_ & new_n420_;
  assign new_n458_ = new_n369_ & new_n423_;
  assign new_n459_ = new_n369_ & new_n421_;
  assign new_n460_ = ~pi31 | ~new_n431_;
  assign new_n461_ = ~pi30 | ~new_n435_;
  assign new_n462_ = ~pi29 | ~new_n439_;
  assign new_n463_ = ~pi28 | ~new_n443_;
  assign new_n464_ = ~pi27 | ~new_n430_;
  assign new_n465_ = ~pi26 | ~new_n434_;
  assign new_n466_ = ~pi25 | ~new_n438_;
  assign new_n467_ = ~pi24 | ~new_n442_;
  assign new_n468_ = ~pi23 | ~new_n429_;
  assign new_n469_ = ~pi22 | ~new_n433_;
  assign new_n470_ = ~pi21 | ~new_n437_;
  assign new_n471_ = ~pi20 | ~new_n441_;
  assign new_n472_ = ~pi19 | ~new_n428_;
  assign new_n473_ = ~pi18 | ~new_n432_;
  assign new_n474_ = ~pi17 | ~new_n436_;
  assign new_n475_ = ~pi16 | ~new_n440_;
  assign new_n476_ = ~pi15 | ~new_n447_;
  assign new_n477_ = ~pi14 | ~new_n451_;
  assign new_n478_ = ~pi13 | ~new_n455_;
  assign new_n479_ = ~pi12 | ~new_n459_;
  assign new_n480_ = ~pi11 | ~new_n446_;
  assign new_n481_ = ~pi10 | ~new_n450_;
  assign new_n482_ = ~pi09 | ~new_n454_;
  assign new_n483_ = ~pi08 | ~new_n458_;
  assign new_n484_ = ~pi07 | ~new_n445_;
  assign new_n485_ = ~pi06 | ~new_n449_;
  assign new_n486_ = ~pi05 | ~new_n453_;
  assign new_n487_ = ~pi04 | ~new_n457_;
  assign new_n488_ = ~pi03 | ~new_n444_;
  assign new_n489_ = ~pi02 | ~new_n448_;
  assign new_n490_ = ~pi01 | ~new_n452_;
  assign new_n491_ = ~pi00 | ~new_n456_;
  assign new_n492_ = ~new_n428_ | ~new_n472_;
  assign new_n493_ = ~new_n429_ | ~new_n468_;
  assign new_n494_ = ~new_n430_ | ~new_n464_;
  assign new_n495_ = ~new_n431_ | ~new_n460_;
  assign new_n496_ = ~new_n432_ | ~new_n473_;
  assign new_n497_ = ~new_n433_ | ~new_n469_;
  assign new_n498_ = ~new_n434_ | ~new_n465_;
  assign new_n499_ = ~new_n435_ | ~new_n461_;
  assign new_n500_ = ~new_n436_ | ~new_n474_;
  assign new_n501_ = ~new_n437_ | ~new_n470_;
  assign new_n502_ = ~new_n438_ | ~new_n466_;
  assign new_n503_ = ~new_n439_ | ~new_n462_;
  assign new_n504_ = ~new_n440_ | ~new_n475_;
  assign new_n505_ = ~new_n441_ | ~new_n471_;
  assign new_n506_ = ~new_n442_ | ~new_n467_;
  assign new_n507_ = ~new_n443_ | ~new_n463_;
  assign new_n508_ = ~new_n444_ | ~new_n488_;
  assign new_n509_ = ~new_n445_ | ~new_n484_;
  assign new_n510_ = ~new_n446_ | ~new_n480_;
  assign new_n511_ = ~new_n447_ | ~new_n476_;
  assign new_n512_ = ~new_n448_ | ~new_n489_;
  assign new_n513_ = ~new_n449_ | ~new_n485_;
  assign new_n514_ = ~new_n450_ | ~new_n481_;
  assign new_n515_ = ~new_n451_ | ~new_n477_;
  assign new_n516_ = ~new_n452_ | ~new_n490_;
  assign new_n517_ = ~new_n453_ | ~new_n486_;
  assign new_n518_ = ~new_n454_ | ~new_n482_;
  assign new_n519_ = ~new_n455_ | ~new_n478_;
  assign new_n520_ = ~new_n456_ | ~new_n491_;
  assign new_n521_ = ~new_n457_ | ~new_n487_;
  assign new_n522_ = ~new_n458_ | ~new_n483_;
  assign new_n523_ = ~new_n459_ | ~new_n479_;
  assign new_n524_ = ~pi31 | ~new_n460_;
  assign new_n525_ = ~pi30 | ~new_n461_;
  assign new_n526_ = ~pi29 | ~new_n462_;
  assign new_n527_ = ~pi28 | ~new_n463_;
  assign new_n528_ = ~pi27 | ~new_n464_;
  assign new_n529_ = ~pi26 | ~new_n465_;
  assign new_n530_ = ~pi25 | ~new_n466_;
  assign new_n531_ = ~pi24 | ~new_n467_;
  assign new_n532_ = ~pi23 | ~new_n468_;
  assign new_n533_ = ~pi22 | ~new_n469_;
  assign new_n534_ = ~pi21 | ~new_n470_;
  assign new_n535_ = ~pi20 | ~new_n471_;
  assign new_n536_ = ~pi19 | ~new_n472_;
  assign new_n537_ = ~pi18 | ~new_n473_;
  assign new_n538_ = ~pi17 | ~new_n474_;
  assign new_n539_ = ~pi16 | ~new_n475_;
  assign new_n540_ = ~pi15 | ~new_n476_;
  assign new_n541_ = ~pi14 | ~new_n477_;
  assign new_n542_ = ~pi13 | ~new_n478_;
  assign new_n543_ = ~pi12 | ~new_n479_;
  assign new_n544_ = ~pi11 | ~new_n480_;
  assign new_n545_ = ~pi10 | ~new_n481_;
  assign new_n546_ = ~pi09 | ~new_n482_;
  assign new_n547_ = ~pi08 | ~new_n483_;
  assign new_n548_ = ~pi07 | ~new_n484_;
  assign new_n549_ = ~pi06 | ~new_n485_;
  assign new_n550_ = ~pi05 | ~new_n486_;
  assign new_n551_ = ~pi04 | ~new_n487_;
  assign new_n552_ = ~pi03 | ~new_n488_;
  assign new_n553_ = ~pi02 | ~new_n489_;
  assign new_n554_ = ~pi01 | ~new_n490_;
  assign new_n555_ = ~pi00 | ~new_n491_;
  assign new_n556_ = ~new_n536_ | ~new_n492_;
  assign new_n557_ = ~new_n532_ | ~new_n493_;
  assign new_n558_ = ~new_n528_ | ~new_n494_;
  assign new_n559_ = ~new_n524_ | ~new_n495_;
  assign new_n560_ = ~new_n537_ | ~new_n496_;
  assign new_n561_ = ~new_n533_ | ~new_n497_;
  assign new_n562_ = ~new_n529_ | ~new_n498_;
  assign new_n563_ = ~new_n525_ | ~new_n499_;
  assign new_n564_ = ~new_n538_ | ~new_n500_;
  assign new_n565_ = ~new_n534_ | ~new_n501_;
  assign new_n566_ = ~new_n530_ | ~new_n502_;
  assign new_n567_ = ~new_n526_ | ~new_n503_;
  assign new_n568_ = ~new_n539_ | ~new_n504_;
  assign new_n569_ = ~new_n535_ | ~new_n505_;
  assign new_n570_ = ~new_n531_ | ~new_n506_;
  assign new_n571_ = ~new_n527_ | ~new_n507_;
  assign new_n572_ = ~new_n552_ | ~new_n508_;
  assign new_n573_ = ~new_n548_ | ~new_n509_;
  assign new_n574_ = ~new_n544_ | ~new_n510_;
  assign new_n575_ = ~new_n540_ | ~new_n511_;
  assign new_n576_ = ~new_n553_ | ~new_n512_;
  assign new_n577_ = ~new_n549_ | ~new_n513_;
  assign new_n578_ = ~new_n545_ | ~new_n514_;
  assign new_n579_ = ~new_n541_ | ~new_n515_;
  assign new_n580_ = ~new_n554_ | ~new_n516_;
  assign new_n581_ = ~new_n550_ | ~new_n517_;
  assign new_n582_ = ~new_n546_ | ~new_n518_;
  assign new_n583_ = ~new_n542_ | ~new_n519_;
  assign new_n584_ = ~new_n555_ | ~new_n520_;
  assign new_n585_ = ~new_n551_ | ~new_n521_;
  assign new_n586_ = ~new_n547_ | ~new_n522_;
  assign new_n587_ = ~new_n543_ | ~new_n523_;
  assign po19 = new_n556_;
  assign po23 = new_n557_;
  assign po27 = new_n558_;
  assign po31 = new_n559_;
  assign po18 = new_n560_;
  assign po22 = new_n561_;
  assign po26 = new_n562_;
  assign po30 = new_n563_;
  assign po17 = new_n564_;
  assign po21 = new_n565_;
  assign po25 = new_n566_;
  assign po29 = new_n567_;
  assign po16 = new_n568_;
  assign po20 = new_n569_;
  assign po24 = new_n570_;
  assign po28 = new_n571_;
  assign po03 = new_n572_;
  assign po07 = new_n573_;
  assign po11 = new_n574_;
  assign po15 = new_n575_;
  assign po02 = new_n576_;
  assign po06 = new_n577_;
  assign po10 = new_n578_;
  assign po14 = new_n579_;
  assign po01 = new_n580_;
  assign po05 = new_n581_;
  assign po09 = new_n582_;
  assign po13 = new_n583_;
  assign po00 = new_n584_;
  assign po04 = new_n585_;
  assign po08 = new_n586_;
  assign po12 = new_n587_;
endmodule


