// Benchmark "pair" written by ABC on Thu Mar 19 13:02:36 2020

module pair ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136;
  wire new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_,
    new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_;
  assign po000 = ~new_n769_;
  assign po001 = ~new_n754_;
  assign po002 = ~new_n739_;
  assign po003 = ~new_n724_;
  assign po004 = ~new_n709_;
  assign po005 = ~new_n1120_;
  assign po006 = ~new_n1105_;
  assign po007 = ~new_n1090_;
  assign po008 = ~new_n1075_;
  assign po009 = ~new_n1060_;
  assign po010 = ~new_n450_ & ~new_n451_;
  assign po011 = ~new_n452_ & ~new_n451_;
  assign po012 = ~new_n453_ & ~new_n451_;
  assign po013 = ~new_n454_ & ~new_n451_;
  assign po014 = ~new_n462_ & ~new_n451_;
  assign po015 = ~new_n463_ & ~new_n451_;
  assign po016 = ~new_n464_ & ~new_n451_;
  assign po017 = ~new_n465_ & ~new_n451_;
  assign po018 = ~new_n467_ & ~new_n451_;
  assign po021 = ~new_n474_ | pi059;
  assign po022 = ~new_n472_ | ~new_n473_;
  assign po023 = ~new_n474_ | ~new_n475_;
  assign po024 = ~new_n493_ | ~new_n494_;
  assign po026 = new_n525_ & ~pi001;
  assign po027 = new_n519_ & ~pi001;
  assign po028 = new_n520_ & ~pi001;
  assign po029 = ~new_n533_;
  assign po030 = ~new_n540_ | ~new_n541_;
  assign po031 = new_n540_ & ~new_n542_;
  assign po032 = new_n540_ & ~new_n543_;
  assign po033 = ~new_n545_ & ~pi001;
  assign po034 = ~new_n552_ & ~pi001;
  assign po035 = ~new_n556_ & ~pi001;
  assign po036 = ~new_n566_ | pi001;
  assign po037 = ~new_n570_ | pi001;
  assign po038 = ~new_n574_ | pi001;
  assign po039 = ~new_n582_ & ~pi001;
  assign po040 = ~new_n586_ | pi001;
  assign po041 = ~new_n590_ | pi001;
  assign po042 = ~pi078 | pi001;
  assign po043 = ~new_n595_ | pi001;
  assign po044 = ~new_n596_ | pi001;
  assign po045 = ~new_n602_ | pi001;
  assign po046 = ~new_n604_ | pi001;
  assign po047 = ~new_n605_ | pi001;
  assign po048 = ~new_n611_ | pi001;
  assign po049 = ~new_n613_ | pi001;
  assign po050 = ~new_n615_ | pi001;
  assign po051 = ~new_n619_ | pi001;
  assign po052 = ~new_n621_ | pi001;
  assign po053 = ~new_n623_ | pi001;
  assign po054 = ~new_n629_ & ~new_n625_ & ~new_n627_ & ~new_n626_;
  assign po055 = ~new_n631_ | pi001;
  assign po056 = (~pi000 & (pi092 | ~new_n442_)) | (pi092 & new_n442_);
  assign po057 = ~new_n632_ & new_n504_;
  assign po058 = ~new_n642_ & new_n504_;
  assign po059 = ~new_n645_ & new_n504_;
  assign po060 = ~new_n650_ | ~new_n651_;
  assign po061 = (new_n482_ & (~new_n504_ | ~new_n652_)) | (new_n504_ & ~new_n652_);
  assign po062 = new_n504_ & ~new_n653_;
  assign po063 = ~new_n663_ & new_n504_;
  assign po064 = ~new_n666_ & new_n504_;
  assign po065 = ~new_n669_ & new_n504_;
  assign po066 = ~new_n677_ | ~new_n678_;
  assign po067 = ~new_n682_ | ~new_n683_;
  assign po068 = ~new_n687_ | ~new_n688_;
  assign po069 = ~new_n697_ & new_n504_;
  assign po070 = ~new_n701_ | ~new_n702_;
  assign po071 = ~new_n706_ | ~new_n707_;
  assign po072 = ~new_n784_ & new_n1025_;
  assign po073 = ~new_n796_ & new_n1025_;
  assign po074 = ~new_n799_ & new_n1025_;
  assign po075 = ~new_n804_ | ~new_n805_;
  assign po076 = (~new_n806_ & new_n1025_) | (new_n999_ & (~new_n806_ | ~new_n1025_));
  assign po077 = new_n1025_ & ~new_n807_;
  assign po078 = ~new_n817_ & new_n1025_;
  assign po079 = ~new_n820_ & new_n1025_;
  assign po080 = ~new_n823_ & new_n1025_;
  assign po081 = ~new_n832_ | ~new_n833_;
  assign po082 = ~new_n837_ | ~new_n838_;
  assign po083 = ~new_n842_ | ~new_n843_;
  assign po084 = ~new_n854_ & new_n1025_;
  assign po085 = ~new_n858_ | ~new_n859_;
  assign po086 = ~new_n863_ | ~new_n864_;
  assign po087 = ~new_n867_ & ~pi024;
  assign po088 = ~new_n875_ & ~pi024;
  assign po089 = ~new_n879_ & ~pi024;
  assign po090 = ~new_n889_ | pi024;
  assign po091 = ~new_n893_ | pi024;
  assign po092 = ~new_n897_ | pi024;
  assign po093 = ~new_n905_ & ~pi024;
  assign po094 = ~new_n909_ | pi024;
  assign po095 = ~new_n913_ | pi024;
  assign po096 = ~pi132 | pi024;
  assign po097 = ~new_n918_ | pi024;
  assign po098 = ~new_n919_ | pi024;
  assign po099 = ~new_n925_ | pi024;
  assign po100 = ~new_n927_ | pi024;
  assign po101 = ~new_n928_ | pi024;
  assign po102 = ~new_n934_ | pi024;
  assign po103 = ~new_n936_ | pi024;
  assign po104 = ~new_n938_ | pi024;
  assign po105 = ~new_n942_ | pi024;
  assign po106 = ~new_n944_ | pi024;
  assign po107 = ~new_n946_ | pi024;
  assign po108 = ~new_n952_ & ~new_n948_ & ~new_n950_ & ~new_n949_;
  assign po109 = ~new_n954_ | pi024;
  assign po110 = ~new_n962_ & ~new_n963_;
  assign po111 = ~new_n964_ & ~new_n963_;
  assign po112 = ~new_n965_ & ~new_n963_;
  assign po113 = ~new_n966_ & ~new_n963_;
  assign po114 = ~new_n974_ & ~new_n963_;
  assign po115 = ~new_n975_ & ~new_n963_;
  assign po116 = ~new_n976_ & ~new_n963_;
  assign po117 = ~new_n977_ & ~new_n963_;
  assign po118 = ~new_n979_ & ~new_n963_;
  assign po121 = ~new_n986_ | pi159;
  assign po122 = ~new_n984_ | ~new_n985_;
  assign po123 = ~new_n986_ | ~new_n987_;
  assign po124 = ~new_n996_ & new_n998_;
  assign po125 = ~new_n997_ & ~pi024;
  assign po126 = ~new_n1010_ | ~new_n998_;
  assign po128 = ~new_n1021_ & ~new_n1022_;
  assign po129 = ~new_n1023_ & ~new_n1022_;
  assign po130 = new_n1043_ & ~pi024;
  assign po131 = new_n1037_ & ~pi024;
  assign po132 = new_n1038_ & ~pi024;
  assign po133 = ~new_n1051_;
  assign po134 = ~new_n1056_ | ~new_n1057_;
  assign po135 = new_n1056_ & ~new_n1058_;
  assign po136 = new_n1056_ & ~new_n1059_;
  assign new_n442_ = new_n624_ | ~pi060;
  assign new_n443_ = pi057 | po021;
  assign new_n444_ = ~new_n443_ & (new_n526_ | ~pi068);
  assign new_n445_ = ~pi046 | ~pi047 | ~pi048 | ~pi049;
  assign new_n446_ = pi046 & new_n489_;
  assign new_n447_ = ~new_n445_ & new_n489_;
  assign new_n448_ = new_n489_ & pi046 & pi047;
  assign new_n449_ = new_n489_ & pi048 & pi046 & pi047;
  assign new_n450_ = pi046 ^ ~new_n489_;
  assign new_n451_ = ~new_n506_ | ~new_n507_ | pi001 | ~new_n487_;
  assign new_n452_ = pi047 ^ ~new_n446_;
  assign new_n453_ = pi048 ^ ~new_n448_;
  assign new_n454_ = pi049 ^ ~new_n449_;
  assign new_n455_ = ~new_n456_ | ~new_n457_;
  assign new_n456_ = ~new_n445_ & ~new_n458_;
  assign new_n457_ = pi053 & new_n489_;
  assign new_n458_ = ~pi052 | ~pi050 | ~pi051;
  assign new_n459_ = new_n489_ & ~new_n445_ & pi050;
  assign new_n460_ = new_n489_ & ~new_n445_ & ~new_n458_;
  assign new_n461_ = new_n489_ & pi051 & ~new_n445_ & pi050;
  assign new_n462_ = pi050 ^ ~new_n447_;
  assign new_n463_ = pi051 ^ ~new_n459_;
  assign new_n464_ = pi052 ^ ~new_n461_;
  assign new_n465_ = pi053 ^ ~new_n460_;
  assign new_n466_ = new_n455_ | ~pi054;
  assign new_n467_ = ~pi054 ^ ~new_n455_;
  assign new_n468_ = ~new_n487_ | pi001;
  assign new_n469_ = ~new_n468_ & (~pi058 | new_n476_);
  assign new_n470_ = ~new_n468_ & (new_n478_ | ~pi059);
  assign new_n471_ = ~new_n472_ | pi058;
  assign new_n472_ = new_n478_ | ~new_n480_ | ~new_n481_;
  assign new_n473_ = ~new_n469_ | ~pi058;
  assign new_n474_ = ~new_n480_ | new_n476_ | ~new_n481_;
  assign new_n475_ = ~new_n470_ | ~pi059;
  assign new_n476_ = ~pi055 | pi056;
  assign new_n477_ = ~po021 & ~pi057;
  assign new_n478_ = ~pi060 | ~new_n479_;
  assign new_n479_ = ~new_n491_ | ~new_n492_;
  assign new_n480_ = ~pi059 & ~pi058;
  assign new_n481_ = ~new_n476_ ^ ~new_n478_;
  assign new_n482_ = ~pi006 & ~new_n497_;
  assign new_n483_ = ~pi054 & new_n484_ & ~pi047;
  assign new_n484_ = ~pi053 & ~pi052 & new_n486_ & ~pi051;
  assign new_n485_ = ~pi048 & ~pi049;
  assign new_n486_ = new_n485_ & ~pi050;
  assign new_n487_ = ~pi064 | pi063 | ~pi062 | pi001;
  assign new_n488_ = ~new_n624_ | ~new_n487_;
  assign new_n489_ = ~new_n444_ | new_n471_;
  assign new_n490_ = ~pi008 & ~new_n443_;
  assign new_n491_ = ~pi065 | pi061;
  assign new_n492_ = pi065 | pi060;
  assign new_n493_ = pi001 | (pi060 & ~new_n624_) | (~pi060 & new_n624_);
  assign new_n494_ = ~new_n498_ & new_n487_;
  assign new_n495_ = ~pi046 & pi047;
  assign new_n496_ = pi046 & new_n483_;
  assign new_n497_ = ~new_n533_ & ~new_n477_;
  assign new_n498_ = ~pi001 & ~pi064 & pi062 & ~pi063;
  assign new_n499_ = new_n483_ & ~pi046;
  assign new_n500_ = ~new_n498_ & (~new_n496_ | new_n533_);
  assign new_n501_ = (new_n505_ | new_n533_) & (new_n526_ | (~pi046 & pi068));
  assign new_n502_ = ~new_n495_ | ((~new_n486_ | ~pi067) & (~pi068 | ~new_n484_) & (~new_n485_ | ~pi066));
  assign new_n503_ = ~new_n501_ | pi005;
  assign new_n504_ = ~pi001 & ~new_n510_;
  assign new_n505_ = ~new_n499_ | (~new_n471_ & ~new_n443_);
  assign new_n506_ = new_n533_ | ~new_n477_ | new_n471_;
  assign new_n507_ = ~pi046 | ~pi068 | new_n526_;
  assign new_n508_ = ~new_n533_ & ~new_n502_;
  assign new_n509_ = ~new_n508_ & ~pi007;
  assign new_n510_ = ~pi001 & ~pi064 & ~pi062 & pi063;
  assign new_n511_ = ~pi002 & ((pi068 & new_n466_) | (~pi054 & (~pi068 | new_n466_)));
  assign new_n512_ = pi105 & pi107 & pi106;
  assign new_n513_ = ~pi001 & pi064 & pi062 & pi063;
  assign new_n514_ = ~new_n513_ & (new_n526_ | new_n476_ | new_n515_ | ~new_n512_);
  assign new_n515_ = ~new_n690_ & ~new_n691_;
  assign new_n516_ = ~pi001 & pi064 & ~pi062 & ~pi063;
  assign new_n517_ = ~new_n498_ & ~new_n516_ & (new_n526_ | ~new_n515_);
  assign new_n518_ = ~new_n513_ & (~pi064 | ~pi063) & (new_n526_ | ~new_n476_ | new_n515_);
  assign new_n519_ = ~new_n524_ | ~new_n518_;
  assign new_n520_ = ~new_n517_ | ~new_n514_;
  assign new_n521_ = new_n533_ | new_n511_;
  assign new_n522_ = new_n526_ | ~new_n515_;
  assign new_n523_ = ~new_n521_ | ~new_n522_;
  assign new_n524_ = ~new_n516_ & ~new_n523_ & ~new_n510_;
  assign new_n525_ = ~new_n527_ | ~new_n529_ | new_n498_;
  assign new_n526_ = ~new_n530_ | ~new_n531_;
  assign new_n527_ = ~new_n510_ | new_n476_;
  assign new_n528_ = ~new_n512_ | new_n515_ | new_n476_;
  assign new_n529_ = ~new_n528_ | new_n526_;
  assign new_n530_ = pi062 & pi063;
  assign new_n531_ = ~pi064 & ~pi001;
  assign new_n532_ = ~new_n534_ | pi064;
  assign new_n533_ = new_n532_ & ~pi001;
  assign new_n534_ = ~pi062 & ~pi063;
  assign new_n535_ = new_n526_ | ~pi066;
  assign new_n536_ = new_n526_ | ~pi067;
  assign new_n537_ = ~pi004 & ~new_n513_;
  assign new_n538_ = ~pi003 & ~new_n516_;
  assign new_n539_ = (~pi066 & (~pi067 | ~pi068)) | (~pi067 & ~pi068);
  assign new_n540_ = new_n539_ & ~pi001 & (pi066 | pi068 | pi067);
  assign new_n541_ = ((~pi067 | new_n538_) & ((~pi066 & (~pi068 | new_n537_)) | (~pi068 & ~new_n537_))) | (~pi067 & ~new_n538_ & (~pi068 | new_n537_));
  assign new_n542_ = ((~pi068 | new_n538_) & ((~pi066 & (~pi067 | ~new_n537_)) | (~pi067 & new_n537_))) | (~pi068 & ~new_n538_ & (~pi066 | new_n537_));
  assign new_n543_ = ((~pi066 | new_n538_) & ((~pi068 & new_n537_) | (~pi067 & (~pi068 | ~new_n537_)))) | (~pi066 & ~new_n538_ & (~pi067 | new_n537_));
  assign new_n544_ = new_n509_ ^ ~pi069;
  assign new_n545_ = (new_n500_ & ~new_n544_) | (~pi099 & (~new_n500_ | ~new_n544_));
  assign new_n546_ = ~pi069 & ~pi070;
  assign new_n547_ = pi070 & pi069;
  assign new_n548_ = pi010 | (~pi071 & ~pi070 & ~pi069);
  assign new_n549_ = pi010 | (pi071 & pi070 & pi069);
  assign new_n550_ = pi069 ^ ~new_n490_;
  assign new_n551_ = ~new_n553_ ^ ~pi070;
  assign new_n552_ = (new_n500_ & ~new_n551_) | (~pi100 & (~new_n500_ | ~new_n551_));
  assign new_n553_ = ~new_n550_ & ~new_n509_;
  assign new_n554_ = (~new_n546_ & (new_n490_ | ~new_n547_)) | (~new_n490_ & ~new_n547_);
  assign new_n555_ = ~new_n557_ ^ ~pi071;
  assign new_n556_ = (new_n500_ & ~new_n555_) | (~pi101 & (~new_n500_ | ~new_n555_));
  assign new_n557_ = ~new_n554_ & ~new_n509_;
  assign new_n558_ = new_n548_ & ~pi072;
  assign new_n559_ = pi072 & new_n549_;
  assign new_n560_ = ~pi073 & new_n548_ & ~pi072;
  assign new_n561_ = new_n549_ & pi073 & pi072;
  assign new_n562_ = pi010 | (~pi074 & ~pi073 & ~pi072 & new_n548_);
  assign new_n563_ = pi010 | (pi074 & pi073 & pi072 & new_n549_);
  assign new_n564_ = (~new_n548_ & (new_n490_ | ~new_n549_)) | (~new_n490_ & ~new_n549_);
  assign new_n565_ = ~new_n567_ ^ ~pi072;
  assign new_n566_ = (new_n500_ & ~new_n565_) | (~pi102 & (~new_n500_ | ~new_n565_));
  assign new_n567_ = ~new_n564_ & ~new_n509_;
  assign new_n568_ = (~new_n558_ & (new_n490_ | ~new_n559_)) | (~new_n490_ & ~new_n559_);
  assign new_n569_ = ~new_n571_ ^ ~pi073;
  assign new_n570_ = (new_n500_ & ~new_n569_) | (~pi103 & (~new_n500_ | ~new_n569_));
  assign new_n571_ = ~new_n568_ & ~new_n509_;
  assign new_n572_ = (~new_n560_ & (new_n490_ | ~new_n561_)) | (~new_n490_ & ~new_n561_);
  assign new_n573_ = ~new_n575_ ^ ~pi074;
  assign new_n574_ = (new_n500_ & ~new_n573_) | (~pi104 & (~new_n500_ | ~new_n573_));
  assign new_n575_ = ~new_n572_ & ~new_n509_;
  assign new_n576_ = new_n562_ & ~pi075;
  assign new_n577_ = pi075 & new_n563_;
  assign new_n578_ = ~pi076 & new_n562_ & ~pi075;
  assign new_n579_ = new_n563_ & pi076 & pi075;
  assign new_n580_ = (~new_n562_ & (new_n490_ | ~new_n563_)) | (~new_n490_ & ~new_n563_);
  assign new_n581_ = ~new_n583_ ^ ~pi075;
  assign new_n582_ = (new_n500_ & ~new_n581_) | (~pi105 & (~new_n500_ | ~new_n581_));
  assign new_n583_ = ~new_n580_ & ~new_n509_;
  assign new_n584_ = (~new_n576_ & (new_n490_ | ~new_n577_)) | (~new_n490_ & ~new_n577_);
  assign new_n585_ = ~new_n587_ ^ ~pi076;
  assign new_n586_ = (new_n500_ & ~new_n585_) | (~pi106 & (~new_n500_ | ~new_n585_));
  assign new_n587_ = ~new_n584_ & ~new_n509_;
  assign new_n588_ = (~new_n578_ & (new_n490_ | ~new_n579_)) | (~new_n490_ & ~new_n579_);
  assign new_n589_ = ~new_n591_ ^ ~pi077;
  assign new_n590_ = (new_n500_ & ~new_n589_) | (~pi107 & (~new_n500_ | ~new_n589_));
  assign new_n591_ = ~new_n588_ & ~new_n509_;
  assign new_n592_ = ~pi067 | pi011;
  assign new_n593_ = pi079 & pi078;
  assign new_n594_ = ~new_n592_ | (pi080 & pi079 & pi078);
  assign new_n595_ = pi078 ^ ~pi079;
  assign new_n596_ = new_n593_ ^ ~pi080;
  assign new_n597_ = ~pi081 | ~new_n600_;
  assign new_n598_ = ~pi083 | ~new_n594_;
  assign new_n599_ = ~pi011 & ~pi066;
  assign new_n600_ = ~new_n598_ | ~new_n599_;
  assign new_n601_ = ~new_n600_ ^ ~pi081;
  assign new_n602_ = (~pi069 & (new_n488_ | ~new_n601_)) | (~new_n488_ & ~new_n601_);
  assign new_n603_ = new_n597_ ^ ~pi082;
  assign new_n604_ = (~pi070 & (new_n488_ | ~new_n603_)) | (~new_n488_ & ~new_n603_);
  assign new_n605_ = new_n594_ ^ ~pi083;
  assign new_n606_ = ~new_n597_ & pi084 & pi082;
  assign new_n607_ = pi082 & ~new_n597_;
  assign new_n608_ = pi085 & new_n606_;
  assign new_n609_ = pi011 | (pi086 & pi085 & new_n606_);
  assign new_n610_ = ~new_n607_ ^ ~pi084;
  assign new_n611_ = (~pi071 & (new_n488_ | ~new_n610_)) | (~new_n488_ & ~new_n610_);
  assign new_n612_ = ~new_n606_ ^ ~pi085;
  assign new_n613_ = (~pi072 & (new_n488_ | ~new_n612_)) | (~new_n488_ & ~new_n612_);
  assign new_n614_ = ~new_n608_ ^ ~pi086;
  assign new_n615_ = (~pi073 & (new_n488_ | ~new_n614_)) | (~new_n488_ & ~new_n614_);
  assign new_n616_ = new_n609_ & pi088 & pi087;
  assign new_n617_ = pi087 & new_n609_;
  assign new_n618_ = ~new_n609_ ^ ~pi087;
  assign new_n619_ = (~pi074 & (new_n488_ | ~new_n618_)) | (~new_n488_ & ~new_n618_);
  assign new_n620_ = ~new_n617_ ^ ~pi088;
  assign new_n621_ = (~pi075 & (new_n488_ | ~new_n620_)) | (~new_n488_ & ~new_n620_);
  assign new_n622_ = ~new_n616_ ^ ~pi089;
  assign new_n623_ = (~pi076 & (new_n488_ | ~new_n622_)) | (~new_n488_ & ~new_n622_);
  assign new_n624_ = ~pi090 | ~new_n600_ | ~pi081;
  assign new_n625_ = ~pi084 | ~pi082;
  assign new_n626_ = ~pi085 | ~pi087 | ~pi086;
  assign new_n627_ = ~pi088 | ~pi091 | ~pi089;
  assign new_n628_ = pi089 & new_n616_;
  assign new_n629_ = new_n488_ & ~pi001;
  assign new_n630_ = ~new_n628_ ^ ~pi091;
  assign new_n631_ = (~pi077 & (new_n488_ | ~new_n630_)) | (~new_n488_ & ~new_n630_);
  assign new_n632_ = new_n503_ ^ ~pi093;
  assign new_n633_ = new_n638_ | (~pi094 & ~pi093);
  assign new_n634_ = ~new_n535_ & ~pi009;
  assign new_n635_ = ~new_n634_ & (pi095 | ~new_n633_);
  assign new_n636_ = new_n638_ | (pi094 & pi093);
  assign new_n637_ = ~new_n634_ & (~pi095 | ~new_n636_);
  assign new_n638_ = ~new_n536_ & ~pi009;
  assign new_n639_ = pi009 | (~pi096 & ~new_n635_);
  assign new_n640_ = pi009 | (pi096 & ~new_n637_);
  assign new_n641_ = pi093 ^ ~new_n482_;
  assign new_n642_ = new_n643_ ^ ~pi094;
  assign new_n643_ = ~new_n641_ & new_n503_;
  assign new_n644_ = (~new_n633_ & (new_n482_ | ~new_n636_)) | (~new_n482_ & ~new_n636_);
  assign new_n645_ = new_n646_ ^ ~pi095;
  assign new_n646_ = ~new_n644_ & new_n503_;
  assign new_n647_ = new_n482_ ? ~new_n635_ : ~new_n637_;
  assign new_n648_ = ~new_n647_ | ~new_n503_;
  assign new_n649_ = new_n648_ ^ ~pi096;
  assign new_n650_ = ~new_n504_ | ~new_n649_;
  assign new_n651_ = new_n504_ | new_n482_;
  assign new_n652_ = pi099 | pi100 | pi101 | pi102;
  assign new_n653_ = ~pi099 | ~pi100 | ~pi101 | ~pi102;
  assign new_n654_ = new_n639_ & ~pi099;
  assign new_n655_ = new_n639_ & pi097;
  assign new_n656_ = pi099 & new_n640_;
  assign new_n657_ = new_n640_ & pi098;
  assign new_n658_ = ~pi100 & new_n639_ & ~pi099;
  assign new_n659_ = new_n640_ & pi100 & pi099;
  assign new_n660_ = ~pi101 & ~pi100 & new_n639_ & ~pi099;
  assign new_n661_ = new_n640_ & pi099 & pi101 & pi100;
  assign new_n662_ = (~new_n639_ & (new_n482_ | ~new_n640_)) | (~new_n482_ & ~new_n640_);
  assign new_n663_ = new_n664_ ^ ~pi099;
  assign new_n664_ = ~new_n662_ & new_n503_;
  assign new_n665_ = (~new_n654_ & (new_n482_ | ~new_n656_)) | (~new_n482_ & ~new_n656_);
  assign new_n666_ = new_n667_ ^ ~pi100;
  assign new_n667_ = ~new_n665_ & new_n503_;
  assign new_n668_ = (~new_n658_ & (new_n482_ | ~new_n659_)) | (~new_n482_ & ~new_n659_);
  assign new_n669_ = new_n670_ ^ ~pi101;
  assign new_n670_ = ~new_n668_ & new_n503_;
  assign new_n671_ = pi009 | (~pi103 & new_n655_);
  assign new_n672_ = ~new_n671_ | pi104;
  assign new_n673_ = pi009 | (pi103 & new_n657_);
  assign new_n674_ = ~pi104 | ~new_n673_;
  assign new_n675_ = (~new_n660_ & (new_n482_ | ~new_n661_)) | (~new_n482_ & ~new_n661_);
  assign new_n676_ = ~new_n679_ ^ ~pi102;
  assign new_n677_ = ~new_n504_ | ~new_n676_;
  assign new_n678_ = new_n504_ | new_n482_;
  assign new_n679_ = ~new_n675_ & new_n503_;
  assign new_n680_ = (~new_n655_ & (new_n482_ | ~new_n657_)) | (~new_n482_ & ~new_n657_);
  assign new_n681_ = ~new_n684_ ^ ~pi103;
  assign new_n682_ = ~new_n504_ | ~new_n681_;
  assign new_n683_ = new_n504_ | new_n482_;
  assign new_n684_ = ~new_n680_ & new_n503_;
  assign new_n685_ = (~new_n671_ & (new_n482_ | ~new_n673_)) | (~new_n482_ & ~new_n673_);
  assign new_n686_ = ~new_n689_ ^ ~pi104;
  assign new_n687_ = ~new_n504_ | ~new_n686_;
  assign new_n688_ = new_n504_ | new_n482_;
  assign new_n689_ = ~new_n685_ & new_n503_;
  assign new_n690_ = pi103 | ~pi101 | pi102;
  assign new_n691_ = pi104 | pi105 | pi106 | pi107;
  assign new_n692_ = ~new_n672_ & ~pi105;
  assign new_n693_ = pi105 & ~new_n674_;
  assign new_n694_ = ~pi106 & ~new_n672_ & ~pi105;
  assign new_n695_ = ~new_n674_ & pi106 & pi105;
  assign new_n696_ = (~new_n482_ & new_n674_) | (new_n672_ & (new_n482_ | new_n674_));
  assign new_n697_ = new_n698_ ^ ~pi105;
  assign new_n698_ = ~new_n696_ & new_n503_;
  assign new_n699_ = (~new_n692_ & (new_n482_ | ~new_n693_)) | (~new_n482_ & ~new_n693_);
  assign new_n700_ = ~new_n703_ ^ ~pi106;
  assign new_n701_ = ~new_n504_ | ~new_n700_;
  assign new_n702_ = new_n504_ | new_n482_;
  assign new_n703_ = ~new_n699_ & new_n503_;
  assign new_n704_ = (~new_n694_ & (new_n482_ | ~new_n695_)) | (~new_n482_ & ~new_n695_);
  assign new_n705_ = ~new_n708_ ^ ~pi107;
  assign new_n706_ = ~new_n504_ | ~new_n705_;
  assign new_n707_ = new_n504_ | new_n482_;
  assign new_n708_ = ~new_n704_ & new_n503_;
  assign new_n709_ = ~new_n721_ & ~new_n722_ & ~new_n723_;
  assign new_n710_ = ~pi022 | ~pi062;
  assign new_n711_ = ~pi021 | ~pi050;
  assign new_n712_ = ~pi020 | new_n503_;
  assign new_n713_ = ~pi019 | ~pi081;
  assign new_n714_ = ~pi018 | new_n624_;
  assign new_n715_ = ~pi017 | ~pi064;
  assign new_n716_ = ~pi016 | new_n504_;
  assign new_n717_ = ~pi015 | ~pi067;
  assign new_n718_ = ~pi014 | ~new_n512_;
  assign new_n719_ = ~pi013 | ~pi099;
  assign new_n720_ = ~pi012 | ~new_n515_;
  assign new_n721_ = ~new_n720_ | ~new_n718_ | ~new_n719_;
  assign new_n722_ = ~new_n710_ | ~new_n711_ | ~new_n712_ | ~new_n713_;
  assign new_n723_ = ~new_n714_ | ~new_n715_ | ~new_n716_ | ~new_n717_;
  assign new_n724_ = ~new_n736_ & ~new_n737_ & ~new_n738_;
  assign new_n725_ = ~pi022 | ~pi046;
  assign new_n726_ = ~pi021 | ~pi051;
  assign new_n727_ = ~pi020 | ~pi078;
  assign new_n728_ = ~pi019 | ~pi082;
  assign new_n729_ = ~pi018 | ~pi087;
  assign new_n730_ = ~pi017 | ~pi063;
  assign new_n731_ = ~pi016 | ~pi068;
  assign new_n732_ = ~pi015 | ~pi066;
  assign new_n733_ = ~pi014 | ~pi093;
  assign new_n734_ = ~pi013 | ~pi100;
  assign new_n735_ = ~pi012 | ~pi104;
  assign new_n736_ = ~new_n735_ | ~new_n733_ | ~new_n734_;
  assign new_n737_ = ~new_n725_ | ~new_n726_ | ~new_n727_ | ~new_n728_;
  assign new_n738_ = ~new_n729_ | ~new_n730_ | ~new_n731_ | ~new_n732_;
  assign new_n739_ = ~new_n751_ & ~new_n752_ & ~new_n753_;
  assign new_n740_ = ~pi022 | ~pi047;
  assign new_n741_ = ~pi021 | ~pi052;
  assign new_n742_ = ~pi020 | ~pi079;
  assign new_n743_ = ~pi019 | ~pi084;
  assign new_n744_ = ~pi018 | ~pi088;
  assign new_n745_ = ~pi017 | ~pi069;
  assign new_n746_ = ~pi016 | ~pi072;
  assign new_n747_ = ~pi015 | ~pi075;
  assign new_n748_ = ~pi014 | ~pi094;
  assign new_n749_ = ~pi013 | ~pi101;
  assign new_n750_ = ~pi012 | ~pi105;
  assign new_n751_ = ~new_n750_ | ~new_n748_ | ~new_n749_;
  assign new_n752_ = ~new_n740_ | ~new_n741_ | ~new_n742_ | ~new_n743_;
  assign new_n753_ = ~new_n744_ | ~new_n745_ | ~new_n746_ | ~new_n747_;
  assign new_n754_ = ~new_n766_ & ~new_n767_ & ~new_n768_;
  assign new_n755_ = ~pi022 | ~pi048;
  assign new_n756_ = ~pi021 | ~pi053;
  assign new_n757_ = ~pi020 | ~pi080;
  assign new_n758_ = ~pi019 | ~pi085;
  assign new_n759_ = ~pi018 | ~pi089;
  assign new_n760_ = ~pi017 | ~pi070;
  assign new_n761_ = ~pi016 | ~pi073;
  assign new_n762_ = ~pi015 | ~pi076;
  assign new_n763_ = ~pi014 | ~pi095;
  assign new_n764_ = ~pi013 | ~pi102;
  assign new_n765_ = ~pi012 | ~pi106;
  assign new_n766_ = ~new_n765_ | ~new_n763_ | ~new_n764_;
  assign new_n767_ = ~new_n755_ | ~new_n756_ | ~new_n757_ | ~new_n758_;
  assign new_n768_ = ~new_n759_ | ~new_n760_ | ~new_n761_ | ~new_n762_;
  assign new_n769_ = ~new_n781_ & ~new_n782_ & ~new_n783_;
  assign new_n770_ = ~pi022 | ~pi049;
  assign new_n771_ = ~pi021 | ~pi054;
  assign new_n772_ = ~pi020 | ~pi083;
  assign new_n773_ = ~pi019 | ~pi086;
  assign new_n774_ = ~pi018 | ~pi091;
  assign new_n775_ = ~pi017 | ~pi071;
  assign new_n776_ = ~pi016 | ~pi074;
  assign new_n777_ = ~pi015 | ~pi077;
  assign new_n778_ = ~pi014 | ~pi096;
  assign new_n779_ = ~pi013 | ~pi103;
  assign new_n780_ = ~pi012 | ~pi107;
  assign new_n781_ = ~new_n780_ | ~new_n778_ | ~new_n779_;
  assign new_n782_ = ~new_n770_ | ~new_n771_ | ~new_n772_ | ~new_n773_;
  assign new_n783_ = ~new_n774_ | ~new_n775_ | ~new_n776_ | ~new_n777_;
  assign new_n784_ = new_n1024_ ^ ~pi108;
  assign new_n785_ = new_n790_ | (~pi109 & ~pi108);
  assign new_n786_ = ~new_n792_ & ~pi032;
  assign new_n787_ = ~new_n786_ & (pi110 | ~new_n785_);
  assign new_n788_ = new_n790_ | (pi109 & pi108);
  assign new_n789_ = ~new_n786_ & (~pi110 | ~new_n788_);
  assign new_n790_ = ~new_n791_ & ~pi032;
  assign new_n791_ = new_n1044_ | ~pi171;
  assign new_n792_ = new_n1044_ | ~pi170;
  assign new_n793_ = pi032 | (~pi111 & ~new_n787_);
  assign new_n794_ = pi032 | (pi111 & ~new_n789_);
  assign new_n795_ = pi108 ^ ~new_n999_;
  assign new_n796_ = new_n797_ ^ ~pi109;
  assign new_n797_ = ~new_n795_ & new_n1024_;
  assign new_n798_ = (~new_n788_ & ~new_n999_) | (~new_n785_ & (~new_n788_ | new_n999_));
  assign new_n799_ = new_n800_ ^ ~pi110;
  assign new_n800_ = ~new_n798_ & new_n1024_;
  assign new_n801_ = new_n999_ ? ~new_n787_ : ~new_n789_;
  assign new_n802_ = ~new_n801_ | ~new_n1024_;
  assign new_n803_ = new_n802_ ^ ~pi111;
  assign new_n804_ = ~new_n1025_ | ~new_n803_;
  assign new_n805_ = new_n1025_ | new_n999_;
  assign new_n806_ = pi114 | pi115 | pi116 | pi117;
  assign new_n807_ = ~pi114 | ~pi115 | ~pi116 | ~pi117;
  assign new_n808_ = new_n793_ & ~pi114;
  assign new_n809_ = new_n793_ & pi112;
  assign new_n810_ = pi114 & new_n794_;
  assign new_n811_ = new_n794_ & pi113;
  assign new_n812_ = ~pi115 & new_n793_ & ~pi114;
  assign new_n813_ = new_n794_ & pi115 & pi114;
  assign new_n814_ = ~pi116 & ~pi115 & new_n793_ & ~pi114;
  assign new_n815_ = new_n794_ & pi114 & pi116 & pi115;
  assign new_n816_ = (~new_n794_ & ~new_n999_) | (~new_n793_ & (~new_n794_ | new_n999_));
  assign new_n817_ = new_n818_ ^ ~pi114;
  assign new_n818_ = ~new_n816_ & new_n1024_;
  assign new_n819_ = (~new_n810_ & ~new_n999_) | (~new_n808_ & (~new_n810_ | new_n999_));
  assign new_n820_ = new_n821_ ^ ~pi115;
  assign new_n821_ = ~new_n819_ & new_n1024_;
  assign new_n822_ = (~new_n813_ & ~new_n999_) | (~new_n812_ & (~new_n813_ | new_n999_));
  assign new_n823_ = new_n824_ ^ ~pi116;
  assign new_n824_ = ~new_n822_ & new_n1024_;
  assign new_n825_ = pi032 | (~pi118 & new_n809_);
  assign new_n826_ = ~new_n825_ | pi119;
  assign new_n827_ = pi032 | (pi118 & new_n811_);
  assign new_n828_ = ~pi119 | ~new_n827_;
  assign new_n829_ = ~pi119 | ~pi118;
  assign new_n830_ = (~new_n815_ & ~new_n999_) | (~new_n814_ & (~new_n815_ | new_n999_));
  assign new_n831_ = ~new_n834_ ^ ~pi117;
  assign new_n832_ = ~new_n1025_ | ~new_n831_;
  assign new_n833_ = new_n1025_ | new_n999_;
  assign new_n834_ = ~new_n830_ & new_n1024_;
  assign new_n835_ = (~new_n811_ & ~new_n999_) | (~new_n809_ & (~new_n811_ | new_n999_));
  assign new_n836_ = ~new_n839_ ^ ~pi118;
  assign new_n837_ = ~new_n1025_ | ~new_n836_;
  assign new_n838_ = new_n1025_ | new_n999_;
  assign new_n839_ = ~new_n835_ & new_n1024_;
  assign new_n840_ = (~new_n827_ & ~new_n999_) | (~new_n825_ & (~new_n827_ | new_n999_));
  assign new_n841_ = ~new_n844_ ^ ~pi119;
  assign new_n842_ = ~new_n1025_ | ~new_n841_;
  assign new_n843_ = new_n1025_ | new_n999_;
  assign new_n844_ = ~new_n840_ & new_n1024_;
  assign new_n845_ = pi118 | ~pi116 | pi117;
  assign new_n846_ = pi119 | pi120 | pi121 | pi122;
  assign new_n847_ = ~new_n826_ & ~pi120;
  assign new_n848_ = pi120 & ~new_n828_;
  assign new_n849_ = ~new_n845_ & ~new_n846_;
  assign new_n850_ = ~pi121 & ~new_n826_ & ~pi120;
  assign new_n851_ = ~new_n828_ & pi121 & pi120;
  assign new_n852_ = ~new_n829_ & pi120 & pi122 & pi121;
  assign new_n853_ = (new_n828_ & ~new_n999_) | (new_n826_ & (new_n828_ | new_n999_));
  assign new_n854_ = new_n855_ ^ ~pi120;
  assign new_n855_ = ~new_n853_ & new_n1024_;
  assign new_n856_ = (~new_n848_ & ~new_n999_) | (~new_n847_ & (~new_n848_ | new_n999_));
  assign new_n857_ = ~new_n860_ ^ ~pi121;
  assign new_n858_ = ~new_n1025_ | ~new_n857_;
  assign new_n859_ = new_n1025_ | new_n999_;
  assign new_n860_ = ~new_n856_ & new_n1024_;
  assign new_n861_ = (~new_n851_ & ~new_n999_) | (~new_n850_ & (~new_n851_ | new_n999_));
  assign new_n862_ = ~new_n865_ ^ ~pi122;
  assign new_n863_ = ~new_n1025_ | ~new_n862_;
  assign new_n864_ = new_n1025_ | new_n999_;
  assign new_n865_ = ~new_n861_ & new_n1024_;
  assign new_n866_ = new_n868_ ^ ~pi123;
  assign new_n867_ = (~new_n866_ & new_n1016_) | (~pi114 & (~new_n866_ | ~new_n1016_));
  assign new_n868_ = ~new_n1029_ & ~pi030;
  assign new_n869_ = ~pi123 & ~pi124;
  assign new_n870_ = pi124 & pi123;
  assign new_n871_ = pi033 | (~pi125 & ~pi124 & ~pi123);
  assign new_n872_ = pi033 | (pi125 & pi124 & pi123);
  assign new_n873_ = pi123 ^ ~new_n1007_;
  assign new_n874_ = ~new_n876_ ^ ~pi124;
  assign new_n875_ = (~new_n874_ & new_n1016_) | (~pi115 & (~new_n874_ | ~new_n1016_));
  assign new_n876_ = ~new_n873_ & ~new_n868_;
  assign new_n877_ = (~new_n870_ & ~new_n1007_) | (~new_n869_ & (~new_n870_ | new_n1007_));
  assign new_n878_ = ~new_n880_ ^ ~pi125;
  assign new_n879_ = (~new_n878_ & new_n1016_) | (~pi116 & (~new_n878_ | ~new_n1016_));
  assign new_n880_ = ~new_n877_ & ~new_n868_;
  assign new_n881_ = new_n871_ & ~pi126;
  assign new_n882_ = pi126 & new_n872_;
  assign new_n883_ = ~pi127 & new_n871_ & ~pi126;
  assign new_n884_ = new_n872_ & pi127 & pi126;
  assign new_n885_ = pi033 | (~pi128 & ~pi127 & ~pi126 & new_n871_);
  assign new_n886_ = pi033 | (pi128 & pi127 & pi126 & new_n872_);
  assign new_n887_ = (~new_n872_ & ~new_n1007_) | (~new_n871_ & (~new_n872_ | new_n1007_));
  assign new_n888_ = ~new_n890_ ^ ~pi126;
  assign new_n889_ = (~new_n888_ & new_n1016_) | (~pi117 & (~new_n888_ | ~new_n1016_));
  assign new_n890_ = ~new_n887_ & ~new_n868_;
  assign new_n891_ = (~new_n882_ & ~new_n1007_) | (~new_n881_ & (~new_n882_ | new_n1007_));
  assign new_n892_ = ~new_n894_ ^ ~pi127;
  assign new_n893_ = (~new_n892_ & new_n1016_) | (~pi118 & (~new_n892_ | ~new_n1016_));
  assign new_n894_ = ~new_n891_ & ~new_n868_;
  assign new_n895_ = (~new_n884_ & ~new_n1007_) | (~new_n883_ & (~new_n884_ | new_n1007_));
  assign new_n896_ = ~new_n898_ ^ ~pi128;
  assign new_n897_ = (~new_n896_ & new_n1016_) | (~pi119 & (~new_n896_ | ~new_n1016_));
  assign new_n898_ = ~new_n895_ & ~new_n868_;
  assign new_n899_ = new_n885_ & ~pi129;
  assign new_n900_ = pi129 & new_n886_;
  assign new_n901_ = ~pi130 & new_n885_ & ~pi129;
  assign new_n902_ = new_n886_ & pi130 & pi129;
  assign new_n903_ = (~new_n886_ & ~new_n1007_) | (~new_n885_ & (~new_n886_ | new_n1007_));
  assign new_n904_ = ~new_n906_ ^ ~pi129;
  assign new_n905_ = (~new_n904_ & new_n1016_) | (~pi120 & (~new_n904_ | ~new_n1016_));
  assign new_n906_ = ~new_n903_ & ~new_n868_;
  assign new_n907_ = (~new_n900_ & ~new_n1007_) | (~new_n899_ & (~new_n900_ | new_n1007_));
  assign new_n908_ = ~new_n910_ ^ ~pi130;
  assign new_n909_ = (~new_n908_ & new_n1016_) | (~pi121 & (~new_n908_ | ~new_n1016_));
  assign new_n910_ = ~new_n907_ & ~new_n868_;
  assign new_n911_ = (~new_n902_ & ~new_n1007_) | (~new_n901_ & (~new_n902_ | new_n1007_));
  assign new_n912_ = ~new_n914_ ^ ~pi131;
  assign new_n913_ = (~new_n912_ & new_n1016_) | (~pi122 & (~new_n912_ | ~new_n1016_));
  assign new_n914_ = ~new_n911_ & ~new_n868_;
  assign new_n915_ = ~pi171 | pi034;
  assign new_n916_ = pi133 & pi132;
  assign new_n917_ = ~new_n915_ | (pi134 & pi133 & pi132);
  assign new_n918_ = pi132 ^ ~pi133;
  assign new_n919_ = new_n916_ ^ ~pi134;
  assign new_n920_ = ~pi135 | ~new_n923_;
  assign new_n921_ = ~pi137 | ~new_n917_;
  assign new_n922_ = ~pi034 & ~pi170;
  assign new_n923_ = ~new_n921_ | ~new_n922_;
  assign new_n924_ = ~new_n923_ ^ ~pi135;
  assign new_n925_ = (~new_n924_ & ~new_n1005_) | (~pi123 & (~new_n924_ | new_n1005_));
  assign new_n926_ = new_n920_ ^ ~pi136;
  assign new_n927_ = (~new_n926_ & ~new_n1005_) | (~pi124 & (~new_n926_ | new_n1005_));
  assign new_n928_ = new_n917_ ^ ~pi137;
  assign new_n929_ = ~new_n920_ & pi138 & pi136;
  assign new_n930_ = pi136 & ~new_n920_;
  assign new_n931_ = pi139 & new_n929_;
  assign new_n932_ = pi034 | (pi140 & pi139 & new_n929_);
  assign new_n933_ = ~new_n930_ ^ ~pi138;
  assign new_n934_ = (~new_n933_ & ~new_n1005_) | (~pi125 & (~new_n933_ | new_n1005_));
  assign new_n935_ = ~new_n929_ ^ ~pi139;
  assign new_n936_ = (~new_n935_ & ~new_n1005_) | (~pi126 & (~new_n935_ | new_n1005_));
  assign new_n937_ = ~new_n931_ ^ ~pi140;
  assign new_n938_ = (~new_n937_ & ~new_n1005_) | (~pi127 & (~new_n937_ | new_n1005_));
  assign new_n939_ = new_n932_ & pi142 & pi141;
  assign new_n940_ = pi141 & new_n932_;
  assign new_n941_ = ~new_n932_ ^ ~pi141;
  assign new_n942_ = (~new_n941_ & ~new_n1005_) | (~pi128 & (~new_n941_ | new_n1005_));
  assign new_n943_ = ~new_n940_ ^ ~pi142;
  assign new_n944_ = (~new_n943_ & ~new_n1005_) | (~pi129 & (~new_n943_ | new_n1005_));
  assign new_n945_ = ~new_n939_ ^ ~pi143;
  assign new_n946_ = (~new_n945_ & ~new_n1005_) | (~pi130 & (~new_n945_ | new_n1005_));
  assign new_n947_ = ~pi144 | ~new_n923_ | ~pi135;
  assign new_n948_ = ~pi138 | ~pi136;
  assign new_n949_ = ~pi139 | ~pi141 | ~pi140;
  assign new_n950_ = ~pi142 | ~pi145 | ~pi143;
  assign new_n951_ = pi143 & new_n939_;
  assign new_n952_ = new_n1005_ & ~pi024;
  assign new_n953_ = ~new_n951_ ^ ~pi145;
  assign new_n954_ = (~new_n953_ & ~new_n1005_) | (~pi131 & (~new_n953_ | new_n1005_));
  assign new_n955_ = pi157 | po121;
  assign new_n956_ = ~new_n955_ & (new_n1044_ | ~pi172);
  assign new_n957_ = ~pi146 | ~pi147 | ~pi148 | ~pi149;
  assign new_n958_ = pi146 & new_n1006_;
  assign new_n959_ = ~new_n957_ & new_n1006_;
  assign new_n960_ = new_n1006_ & pi146 & pi147;
  assign new_n961_ = new_n1006_ & pi148 & pi146 & pi147;
  assign new_n962_ = pi146 ^ ~new_n1006_;
  assign new_n963_ = ~new_n1027_ | ~new_n1028_ | pi024 | ~new_n1004_;
  assign new_n964_ = pi147 ^ ~new_n958_;
  assign new_n965_ = pi148 ^ ~new_n960_;
  assign new_n966_ = pi149 ^ ~new_n961_;
  assign new_n967_ = ~new_n968_ | ~new_n969_;
  assign new_n968_ = ~new_n957_ & ~new_n970_;
  assign new_n969_ = pi153 & new_n1006_;
  assign new_n970_ = ~pi152 | ~pi150 | ~pi151;
  assign new_n971_ = new_n1006_ & ~new_n957_ & pi150;
  assign new_n972_ = new_n1006_ & ~new_n957_ & ~new_n970_;
  assign new_n973_ = new_n1006_ & pi151 & ~new_n957_ & pi150;
  assign new_n974_ = pi150 ^ ~new_n959_;
  assign new_n975_ = pi151 ^ ~new_n971_;
  assign new_n976_ = pi152 ^ ~new_n973_;
  assign new_n977_ = pi153 ^ ~new_n972_;
  assign new_n978_ = new_n967_ | ~pi154;
  assign new_n979_ = ~pi154 ^ ~new_n967_;
  assign new_n980_ = pi024 | ~new_n1004_;
  assign new_n981_ = ~new_n980_ & (~pi158 | new_n988_);
  assign new_n982_ = ~new_n980_ & (new_n990_ | ~pi159);
  assign new_n983_ = ~new_n984_ | pi158;
  assign new_n984_ = new_n990_ | ~new_n992_ | ~new_n993_;
  assign new_n985_ = ~new_n981_ | ~pi158;
  assign new_n986_ = ~new_n992_ | new_n988_ | ~new_n993_;
  assign new_n987_ = ~new_n982_ | ~pi159;
  assign new_n988_ = ~pi155 | pi156;
  assign new_n989_ = ~po121 & ~pi157;
  assign new_n990_ = ~pi161 | ~new_n991_;
  assign new_n991_ = ~new_n1008_ | ~new_n1009_;
  assign new_n992_ = ~pi159 & ~pi158;
  assign new_n993_ = ~new_n988_ ^ ~new_n990_;
  assign new_n994_ = ~po126 | pi162;
  assign new_n995_ = ~pi161 & ~pi160;
  assign new_n996_ = ~pi024 & ((~new_n994_ & ~new_n995_) | (~pi160 & (new_n994_ | ~new_n995_)));
  assign new_n997_ = new_n998_ & ((~pi161 & new_n994_) | (~pi160 & (~pi161 | ~new_n994_)));
  assign new_n998_ = ~new_n1014_ & new_n1004_;
  assign new_n999_ = ~pi029 & ~new_n1013_;
  assign new_n1000_ = ~pi154 & new_n1001_ & ~pi147;
  assign new_n1001_ = ~pi153 & ~pi152 & new_n1003_ & ~pi151;
  assign new_n1002_ = ~pi148 & ~pi149;
  assign new_n1003_ = new_n1002_ & ~pi150;
  assign new_n1004_ = ~pi168 | pi167 | ~pi166 | pi024;
  assign new_n1005_ = ~new_n947_ | ~new_n1004_;
  assign new_n1006_ = ~new_n956_ | new_n983_;
  assign new_n1007_ = ~pi031 & ~new_n955_;
  assign new_n1008_ = ~pi169 | pi163;
  assign new_n1009_ = pi169 | pi161;
  assign new_n1010_ = pi024 | (pi162 & ~new_n947_) | (~pi162 & new_n947_);
  assign new_n1011_ = ~pi146 & pi147;
  assign new_n1012_ = pi146 & new_n1000_;
  assign new_n1013_ = ~new_n1051_ & ~new_n989_;
  assign new_n1014_ = ~pi024 & ~pi168 & pi166 & ~pi167;
  assign new_n1015_ = new_n1000_ & ~pi146;
  assign new_n1016_ = ~new_n1014_ & (~new_n1012_ | new_n1051_);
  assign new_n1017_ = pi165 & ~pi164;
  assign new_n1018_ = (new_n1026_ | new_n1051_) & (~new_n1017_ | (~pi146 & pi172));
  assign new_n1019_ = ~new_n1011_ | ((~pi172 | ~new_n1001_) & (~pi170 | ~new_n1002_) & (~pi171 | ~new_n1003_));
  assign new_n1020_ = ~new_n1044_ & pi164;
  assign new_n1021_ = ~pi164 ^ ~new_n1044_;
  assign new_n1022_ = pi024 | new_n1017_;
  assign new_n1023_ = pi165 ^ ~new_n1020_;
  assign new_n1024_ = ~new_n1018_ | pi028;
  assign new_n1025_ = ~pi024 & ~new_n1030_;
  assign new_n1026_ = ~new_n1015_ | (~new_n983_ & ~new_n955_);
  assign new_n1027_ = new_n1051_ | ~new_n989_ | new_n983_;
  assign new_n1028_ = ~pi146 | ~pi172 | new_n1044_;
  assign new_n1029_ = ~new_n1051_ & ~new_n1019_;
  assign new_n1030_ = ~pi024 & ~pi168 & ~pi166 & pi167;
  assign new_n1031_ = ~pi025 & ((pi172 & new_n978_) | (~pi154 & (~pi172 | new_n978_)));
  assign new_n1032_ = ~pi024 & pi168 & pi166 & pi167;
  assign new_n1033_ = ~new_n1032_ & (new_n1044_ | new_n988_ | new_n849_ | ~new_n852_);
  assign new_n1034_ = ~pi024 & pi168 & ~pi166 & ~pi167;
  assign new_n1035_ = ~new_n1014_ & ~new_n1034_ & (new_n1044_ | ~new_n849_);
  assign new_n1036_ = ~new_n1032_ & (~pi168 | ~pi167) & (new_n1044_ | ~new_n988_ | new_n849_);
  assign new_n1037_ = ~new_n1042_ | ~new_n1036_;
  assign new_n1038_ = ~new_n1035_ | ~new_n1033_;
  assign new_n1039_ = new_n1051_ | new_n1031_;
  assign new_n1040_ = new_n1044_ | ~new_n849_;
  assign new_n1041_ = ~new_n1039_ | ~new_n1040_;
  assign new_n1042_ = ~new_n1034_ & ~new_n1041_ & ~new_n1030_;
  assign new_n1043_ = ~new_n1045_ | ~new_n1047_ | new_n1014_;
  assign new_n1044_ = ~new_n1048_ | ~new_n1049_;
  assign new_n1045_ = ~new_n1030_ | new_n988_;
  assign new_n1046_ = ~new_n852_ | new_n849_ | new_n988_;
  assign new_n1047_ = ~new_n1046_ | new_n1044_;
  assign new_n1048_ = pi166 & pi167;
  assign new_n1049_ = ~pi168 & ~pi024;
  assign new_n1050_ = ~new_n1052_ | pi168;
  assign new_n1051_ = new_n1050_ & ~pi024;
  assign new_n1052_ = ~pi166 & ~pi167;
  assign new_n1053_ = ~pi027 & ~new_n1032_;
  assign new_n1054_ = ~pi026 & ~new_n1034_;
  assign new_n1055_ = (~pi170 & (~pi171 | ~pi172)) | (~pi171 & ~pi172);
  assign new_n1056_ = new_n1055_ & ~pi024 & (pi170 | pi172 | pi171);
  assign new_n1057_ = ((~pi171 | new_n1054_) & ((~pi170 & (~pi172 | new_n1053_)) | (~pi172 & ~new_n1053_))) | (~pi171 & ~new_n1054_ & (~pi172 | new_n1053_));
  assign new_n1058_ = ((~pi172 | new_n1054_) & ((~pi170 & (~pi171 | ~new_n1053_)) | (~pi171 & new_n1053_))) | (~pi172 & ~new_n1054_ & (~pi170 | new_n1053_));
  assign new_n1059_ = ((~pi170 | new_n1054_) & ((~pi172 & new_n1053_) | (~pi171 & (~pi172 | ~new_n1053_)))) | (~pi170 & ~new_n1054_ & (~pi171 | new_n1053_));
  assign new_n1060_ = ~new_n1072_ & ~new_n1073_ & ~new_n1074_;
  assign new_n1061_ = ~pi045 | ~pi166;
  assign new_n1062_ = ~pi044 | ~pi150;
  assign new_n1063_ = ~pi043 | new_n1024_;
  assign new_n1064_ = ~pi042 | ~pi135;
  assign new_n1065_ = ~pi041 | new_n947_;
  assign new_n1066_ = ~pi040 | ~pi168;
  assign new_n1067_ = ~pi039 | new_n1025_;
  assign new_n1068_ = ~pi038 | ~pi171;
  assign new_n1069_ = ~pi037 | ~new_n852_;
  assign new_n1070_ = ~pi036 | ~pi114;
  assign new_n1071_ = ~pi035 | ~new_n849_;
  assign new_n1072_ = ~new_n1071_ | ~new_n1069_ | ~new_n1070_;
  assign new_n1073_ = ~new_n1061_ | ~new_n1062_ | ~new_n1063_ | ~new_n1064_;
  assign new_n1074_ = ~new_n1065_ | ~new_n1066_ | ~new_n1067_ | ~new_n1068_;
  assign new_n1075_ = ~new_n1087_ & ~new_n1088_ & ~new_n1089_;
  assign new_n1076_ = ~pi045 | ~pi146;
  assign new_n1077_ = ~pi044 | ~pi151;
  assign new_n1078_ = ~pi043 | ~pi132;
  assign new_n1079_ = ~pi042 | ~pi136;
  assign new_n1080_ = ~pi041 | ~pi141;
  assign new_n1081_ = ~pi040 | ~pi167;
  assign new_n1082_ = ~pi039 | ~pi172;
  assign new_n1083_ = ~pi038 | ~pi170;
  assign new_n1084_ = ~pi037 | ~pi108;
  assign new_n1085_ = ~pi036 | ~pi115;
  assign new_n1086_ = ~pi035 | ~pi119;
  assign new_n1087_ = ~new_n1086_ | ~new_n1084_ | ~new_n1085_;
  assign new_n1088_ = ~new_n1076_ | ~new_n1077_ | ~new_n1078_ | ~new_n1079_;
  assign new_n1089_ = ~new_n1080_ | ~new_n1081_ | ~new_n1082_ | ~new_n1083_;
  assign new_n1090_ = ~new_n1102_ & ~new_n1103_ & ~new_n1104_;
  assign new_n1091_ = ~pi045 | ~pi147;
  assign new_n1092_ = ~pi044 | ~pi152;
  assign new_n1093_ = ~pi043 | ~pi133;
  assign new_n1094_ = ~pi042 | ~pi138;
  assign new_n1095_ = ~pi041 | ~pi142;
  assign new_n1096_ = ~pi040 | ~pi123;
  assign new_n1097_ = ~pi039 | ~pi126;
  assign new_n1098_ = ~pi038 | ~pi129;
  assign new_n1099_ = ~pi037 | ~pi109;
  assign new_n1100_ = ~pi036 | ~pi116;
  assign new_n1101_ = ~pi035 | ~pi120;
  assign new_n1102_ = ~new_n1101_ | ~new_n1099_ | ~new_n1100_;
  assign new_n1103_ = ~new_n1091_ | ~new_n1092_ | ~new_n1093_ | ~new_n1094_;
  assign new_n1104_ = ~new_n1095_ | ~new_n1096_ | ~new_n1097_ | ~new_n1098_;
  assign new_n1105_ = ~new_n1117_ & ~new_n1118_ & ~new_n1119_;
  assign new_n1106_ = ~pi045 | ~pi148;
  assign new_n1107_ = ~pi044 | ~pi153;
  assign new_n1108_ = ~pi043 | ~pi134;
  assign new_n1109_ = ~pi042 | ~pi139;
  assign new_n1110_ = ~pi041 | ~pi143;
  assign new_n1111_ = ~pi040 | ~pi124;
  assign new_n1112_ = ~pi039 | ~pi127;
  assign new_n1113_ = ~pi038 | ~pi130;
  assign new_n1114_ = ~pi037 | ~pi110;
  assign new_n1115_ = ~pi036 | ~pi117;
  assign new_n1116_ = ~pi035 | ~pi121;
  assign new_n1117_ = ~new_n1116_ | ~new_n1114_ | ~new_n1115_;
  assign new_n1118_ = ~new_n1106_ | ~new_n1107_ | ~new_n1108_ | ~new_n1109_;
  assign new_n1119_ = ~new_n1110_ | ~new_n1111_ | ~new_n1112_ | ~new_n1113_;
  assign new_n1120_ = ~new_n1132_ & ~new_n1133_ & ~new_n1134_;
  assign new_n1121_ = ~pi045 | ~pi149;
  assign new_n1122_ = ~pi044 | ~pi154;
  assign new_n1123_ = ~pi043 | ~pi137;
  assign new_n1124_ = ~pi042 | ~pi140;
  assign new_n1125_ = ~pi041 | ~pi145;
  assign new_n1126_ = ~pi040 | ~pi125;
  assign new_n1127_ = ~pi039 | ~pi128;
  assign new_n1128_ = ~pi038 | ~pi131;
  assign new_n1129_ = ~pi037 | ~pi111;
  assign new_n1130_ = ~pi036 | ~pi118;
  assign new_n1131_ = ~pi035 | ~pi122;
  assign new_n1132_ = ~new_n1131_ | ~new_n1129_ | ~new_n1130_;
  assign new_n1133_ = ~new_n1121_ | ~new_n1122_ | ~new_n1123_ | ~new_n1124_;
  assign new_n1134_ = ~new_n1125_ | ~new_n1126_ | ~new_n1127_ | ~new_n1128_;
  assign po019 = pi000;
  assign po020 = pi055;
  assign po025 = pi060;
  assign po119 = pi023;
  assign po120 = pi155;
  assign po127 = pi161;
endmodule


