// Benchmark "i7" written by ABC on Thu Mar 19 13:02:36 2020

module i7 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47,
    po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46,
    po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58,
    po59, po60, po61, po62, po63, po64, po65, po66;
  wire new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n299_, new_n301_, new_n303_, new_n305_, new_n307_,
    new_n309_, new_n311_, new_n313_, new_n315_, new_n317_, new_n319_,
    new_n321_, new_n323_, new_n325_, new_n327_, new_n329_, new_n331_,
    new_n333_, new_n335_, new_n337_, new_n339_, new_n341_, new_n343_,
    new_n345_, new_n347_, new_n349_, new_n351_, new_n353_, new_n354_,
    new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_,
    new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_,
    new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_,
    new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_,
    new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_,
    new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n445_,
    new_n447_, new_n449_, new_n451_, new_n453_, new_n455_, new_n457_,
    new_n459_, new_n461_, new_n463_, new_n465_, new_n467_, new_n469_,
    new_n471_, new_n473_, new_n475_, new_n477_, new_n479_, new_n481_,
    new_n483_, new_n485_, new_n487_, new_n489_, new_n491_, new_n493_,
    new_n495_, new_n497_, new_n499_, new_n501_, new_n503_, new_n505_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n581_, new_n583_, new_n585_, new_n587_, new_n589_,
    new_n591_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_;
  assign new_n267_ = ~pi000;
  assign new_n268_ = pi002 & pi001 & new_n267_;
  assign new_n269_ = pi002 & pi003 & new_n267_;
  assign new_n270_ = pi002 & pi004 & new_n267_;
  assign new_n271_ = pi002 & pi005 & new_n267_;
  assign new_n272_ = pi002 & pi006 & new_n267_;
  assign new_n273_ = pi002 & pi007 & new_n267_;
  assign new_n274_ = pi002 & pi008 & new_n267_;
  assign new_n275_ = pi002 & pi009 & new_n267_;
  assign new_n276_ = pi002 & pi010 & new_n267_;
  assign new_n277_ = pi002 & pi011 & new_n267_;
  assign new_n278_ = pi002 & pi012 & new_n267_;
  assign new_n279_ = pi002 & pi013 & new_n267_;
  assign new_n280_ = pi002 & pi014 & new_n267_;
  assign new_n281_ = pi002 & pi015 & new_n267_;
  assign new_n282_ = pi002 & pi016 & new_n267_;
  assign new_n283_ = pi002 & pi017 & new_n267_;
  assign new_n284_ = pi002 & pi018 & new_n267_;
  assign new_n285_ = pi002 & pi019 & new_n267_;
  assign new_n286_ = pi002 & pi020 & new_n267_;
  assign new_n287_ = pi002 & pi021 & new_n267_;
  assign new_n288_ = pi002 & pi022 & new_n267_;
  assign new_n289_ = pi002 & pi023 & new_n267_;
  assign new_n290_ = pi002 & pi024 & new_n267_;
  assign new_n291_ = pi002 & pi025 & new_n267_;
  assign new_n292_ = pi002 & pi026 & new_n267_;
  assign new_n293_ = pi002 & pi027 & new_n267_;
  assign new_n294_ = pi002 & pi028 & new_n267_;
  assign new_n295_ = pi002 & pi029 & new_n267_;
  assign new_n296_ = ~pi002;
  assign new_n297_ = new_n296_ & pi030 & new_n267_;
  assign po00 = new_n353_ | new_n381_ | new_n268_ | new_n297_;
  assign new_n299_ = new_n296_ & pi031 & new_n267_;
  assign po01 = new_n354_ | new_n382_ | new_n269_ | new_n299_;
  assign new_n301_ = new_n296_ & pi032 & new_n267_;
  assign po02 = new_n355_ | new_n383_ | new_n270_ | new_n301_;
  assign new_n303_ = new_n296_ & pi033 & new_n267_;
  assign po03 = new_n356_ | new_n384_ | new_n271_ | new_n303_;
  assign new_n305_ = new_n296_ & pi034 & new_n267_;
  assign po04 = new_n357_ | new_n385_ | new_n272_ | new_n305_;
  assign new_n307_ = new_n296_ & pi035 & new_n267_;
  assign po05 = new_n358_ | new_n386_ | new_n273_ | new_n307_;
  assign new_n309_ = new_n296_ & pi036 & new_n267_;
  assign po06 = new_n359_ | new_n387_ | new_n274_ | new_n309_;
  assign new_n311_ = new_n296_ & pi037 & new_n267_;
  assign po07 = new_n360_ | new_n388_ | new_n275_ | new_n311_;
  assign new_n313_ = new_n296_ & pi038 & new_n267_;
  assign po08 = new_n361_ | new_n389_ | new_n276_ | new_n313_;
  assign new_n315_ = new_n296_ & pi039 & new_n267_;
  assign po09 = new_n362_ | new_n390_ | new_n277_ | new_n315_;
  assign new_n317_ = new_n296_ & pi040 & new_n267_;
  assign po10 = new_n363_ | new_n391_ | new_n278_ | new_n317_;
  assign new_n319_ = new_n296_ & pi041 & new_n267_;
  assign po11 = new_n364_ | new_n392_ | new_n279_ | new_n319_;
  assign new_n321_ = new_n296_ & pi042 & new_n267_;
  assign po12 = new_n365_ | new_n393_ | new_n280_ | new_n321_;
  assign new_n323_ = new_n296_ & pi043 & new_n267_;
  assign po13 = new_n366_ | new_n394_ | new_n281_ | new_n323_;
  assign new_n325_ = new_n296_ & pi044 & new_n267_;
  assign po14 = new_n367_ | new_n395_ | new_n282_ | new_n325_;
  assign new_n327_ = new_n296_ & pi045 & new_n267_;
  assign po15 = new_n368_ | new_n396_ | new_n283_ | new_n327_;
  assign new_n329_ = new_n296_ & pi046 & new_n267_;
  assign po16 = new_n369_ | new_n397_ | new_n284_ | new_n329_;
  assign new_n331_ = new_n296_ & pi047 & new_n267_;
  assign po17 = new_n370_ | new_n398_ | new_n285_ | new_n331_;
  assign new_n333_ = new_n296_ & pi048 & new_n267_;
  assign po18 = new_n371_ | new_n399_ | new_n286_ | new_n333_;
  assign new_n335_ = new_n296_ & pi049 & new_n267_;
  assign po19 = new_n372_ | new_n400_ | new_n287_ | new_n335_;
  assign new_n337_ = new_n296_ & pi050 & new_n267_;
  assign po20 = new_n373_ | new_n401_ | new_n288_ | new_n337_;
  assign new_n339_ = new_n296_ & pi051 & new_n267_;
  assign po21 = new_n374_ | new_n402_ | new_n289_ | new_n339_;
  assign new_n341_ = new_n296_ & pi052 & new_n267_;
  assign po22 = new_n375_ | new_n403_ | new_n290_ | new_n341_;
  assign new_n343_ = new_n296_ & pi053 & new_n267_;
  assign po23 = new_n376_ | new_n404_ | new_n291_ | new_n343_;
  assign new_n345_ = new_n296_ & pi054 & new_n267_;
  assign po24 = new_n377_ | new_n405_ | new_n292_ | new_n345_;
  assign new_n347_ = new_n296_ & pi055 & new_n267_;
  assign po25 = new_n378_ | new_n406_ | new_n293_ | new_n347_;
  assign new_n349_ = new_n296_ & pi056 & new_n267_;
  assign po26 = new_n379_ | new_n407_ | new_n294_ | new_n349_;
  assign new_n351_ = new_n296_ & pi057 & new_n267_;
  assign po27 = new_n380_ | new_n408_ | new_n295_ | new_n351_;
  assign new_n353_ = pi002 & pi058 & pi000;
  assign new_n354_ = pi002 & pi059 & pi000;
  assign new_n355_ = pi002 & pi060 & pi000;
  assign new_n356_ = pi002 & pi061 & pi000;
  assign new_n357_ = pi002 & pi062 & pi000;
  assign new_n358_ = pi002 & pi063 & pi000;
  assign new_n359_ = pi002 & pi064 & pi000;
  assign new_n360_ = pi002 & pi065 & pi000;
  assign new_n361_ = pi002 & pi066 & pi000;
  assign new_n362_ = pi002 & pi067 & pi000;
  assign new_n363_ = pi002 & pi068 & pi000;
  assign new_n364_ = pi002 & pi069 & pi000;
  assign new_n365_ = pi002 & pi070 & pi000;
  assign new_n366_ = pi002 & pi071 & pi000;
  assign new_n367_ = pi002 & pi072 & pi000;
  assign new_n368_ = pi002 & pi073 & pi000;
  assign new_n369_ = pi002 & pi074 & pi000;
  assign new_n370_ = pi002 & pi075 & pi000;
  assign new_n371_ = pi002 & pi076 & pi000;
  assign new_n372_ = pi002 & pi077 & pi000;
  assign new_n373_ = pi002 & pi078 & pi000;
  assign new_n374_ = pi002 & pi079 & pi000;
  assign new_n375_ = pi002 & pi080 & pi000;
  assign new_n376_ = pi002 & pi081 & pi000;
  assign new_n377_ = pi002 & pi082 & pi000;
  assign new_n378_ = pi002 & pi083 & pi000;
  assign new_n379_ = pi002 & pi084 & pi000;
  assign new_n380_ = pi002 & pi085 & pi000;
  assign new_n381_ = new_n296_ & new_n634_ & pi000;
  assign new_n382_ = new_n296_ & new_n633_ & pi000;
  assign new_n383_ = new_n296_ & new_n632_ & pi000;
  assign new_n384_ = new_n296_ & new_n631_ & pi000;
  assign new_n385_ = new_n296_ & new_n630_ & pi000;
  assign new_n386_ = new_n296_ & new_n629_ & pi000;
  assign new_n387_ = new_n296_ & new_n628_ & pi000;
  assign new_n388_ = new_n296_ & new_n627_ & pi000;
  assign new_n389_ = new_n296_ & new_n626_ & pi000;
  assign new_n390_ = new_n296_ & new_n625_ & pi000;
  assign new_n391_ = new_n296_ & new_n624_ & pi000;
  assign new_n392_ = new_n296_ & new_n623_ & pi000;
  assign new_n393_ = new_n296_ & new_n622_ & pi000;
  assign new_n394_ = new_n296_ & new_n621_ & pi000;
  assign new_n395_ = new_n296_ & new_n620_ & pi000;
  assign new_n396_ = new_n296_ & new_n619_ & pi000;
  assign new_n397_ = new_n296_ & new_n618_ & pi000;
  assign new_n398_ = new_n296_ & new_n617_ & pi000;
  assign new_n399_ = new_n296_ & new_n616_ & pi000;
  assign new_n400_ = new_n296_ & new_n615_ & pi000;
  assign new_n401_ = new_n296_ & new_n614_ & pi000;
  assign new_n402_ = new_n296_ & new_n613_ & pi000;
  assign new_n403_ = new_n296_ & new_n612_ & pi000;
  assign new_n404_ = new_n296_ & new_n611_ & pi000;
  assign new_n405_ = new_n296_ & new_n610_ & pi000;
  assign new_n406_ = new_n296_ & new_n609_ & pi000;
  assign new_n407_ = new_n296_ & new_n608_ & pi000;
  assign new_n408_ = new_n296_ & new_n607_ & pi000;
  assign new_n409_ = ~pi000;
  assign new_n410_ = pi087 & new_n409_ & pi086 & pi002;
  assign new_n411_ = pi087 & new_n409_ & pi088 & pi002;
  assign new_n412_ = pi087 & new_n409_ & pi089 & pi002;
  assign new_n413_ = pi087 & new_n409_ & pi090 & pi002;
  assign new_n414_ = pi087 & new_n409_ & pi091 & pi002;
  assign new_n415_ = pi087 & new_n409_ & pi092 & pi002;
  assign new_n416_ = pi087 & new_n409_ & pi093 & pi002;
  assign new_n417_ = pi087 & new_n409_ & pi094 & pi002;
  assign new_n418_ = pi087 & new_n409_ & pi095 & pi002;
  assign new_n419_ = pi087 & new_n409_ & pi096 & pi002;
  assign new_n420_ = pi087 & new_n409_ & pi097 & pi002;
  assign new_n421_ = pi087 & new_n409_ & pi098 & pi002;
  assign new_n422_ = pi087 & new_n409_ & pi099 & pi002;
  assign new_n423_ = pi087 & new_n409_ & pi100 & pi002;
  assign new_n424_ = pi087 & new_n409_ & pi101 & pi002;
  assign new_n425_ = pi087 & new_n409_ & pi102 & pi002;
  assign new_n426_ = pi087 & new_n409_ & pi103 & pi002;
  assign new_n427_ = pi087 & new_n409_ & pi104 & pi002;
  assign new_n428_ = pi087 & new_n409_ & pi105 & pi002;
  assign new_n429_ = pi087 & new_n409_ & pi106 & pi002;
  assign new_n430_ = pi087 & new_n409_ & pi107 & pi002;
  assign new_n431_ = pi087 & new_n409_ & pi108 & pi002;
  assign new_n432_ = pi087 & new_n409_ & pi109 & pi002;
  assign new_n433_ = pi087 & new_n409_ & pi110 & pi002;
  assign new_n434_ = pi087 & new_n409_ & pi111 & pi002;
  assign new_n435_ = pi087 & new_n409_ & pi112 & pi002;
  assign new_n436_ = pi087 & new_n409_ & pi113 & pi002;
  assign new_n437_ = pi087 & new_n409_ & pi114 & pi002;
  assign new_n438_ = pi087 & new_n409_ & pi115 & pi002;
  assign new_n439_ = pi087 & new_n409_ & pi116 & pi002;
  assign new_n440_ = pi087 & new_n409_ & pi117 & pi002;
  assign new_n441_ = pi087 & new_n409_ & pi118 & pi002;
  assign new_n442_ = ~pi002;
  assign new_n443_ = pi087 & new_n409_ & pi119 & new_n442_;
  assign po28 = new_n539_ | new_n572_ | new_n507_ | new_n410_ | new_n443_;
  assign new_n445_ = pi087 & new_n409_ & pi120 & new_n442_;
  assign po29 = new_n540_ | new_n572_ | new_n508_ | new_n411_ | new_n445_;
  assign new_n447_ = pi087 & new_n409_ & pi121 & new_n442_;
  assign po30 = new_n541_ | new_n572_ | new_n509_ | new_n412_ | new_n447_;
  assign new_n449_ = pi087 & new_n409_ & pi122 & new_n442_;
  assign po31 = new_n542_ | new_n572_ | new_n510_ | new_n413_ | new_n449_;
  assign new_n451_ = pi087 & new_n409_ & pi123 & new_n442_;
  assign po32 = new_n543_ | new_n572_ | new_n511_ | new_n414_ | new_n451_;
  assign new_n453_ = pi087 & new_n409_ & pi124 & new_n442_;
  assign po33 = new_n544_ | new_n572_ | new_n512_ | new_n415_ | new_n453_;
  assign new_n455_ = pi087 & new_n409_ & pi125 & new_n442_;
  assign po34 = new_n545_ | new_n572_ | new_n513_ | new_n416_ | new_n455_;
  assign new_n457_ = pi087 & new_n409_ & pi126 & new_n442_;
  assign po35 = new_n546_ | new_n572_ | new_n514_ | new_n417_ | new_n457_;
  assign new_n459_ = pi087 & new_n409_ & pi127 & new_n442_;
  assign po36 = new_n547_ | new_n572_ | new_n515_ | new_n418_ | new_n459_;
  assign new_n461_ = pi087 & new_n409_ & pi128 & new_n442_;
  assign po37 = new_n548_ | new_n572_ | new_n516_ | new_n419_ | new_n461_;
  assign new_n463_ = pi087 & new_n409_ & pi129 & new_n442_;
  assign po38 = new_n549_ | new_n572_ | new_n517_ | new_n420_ | new_n463_;
  assign new_n465_ = pi087 & new_n409_ & pi130 & new_n442_;
  assign po39 = new_n550_ | new_n572_ | new_n518_ | new_n421_ | new_n465_;
  assign new_n467_ = pi087 & new_n409_ & pi131 & new_n442_;
  assign po40 = new_n551_ | new_n572_ | new_n519_ | new_n422_ | new_n467_;
  assign new_n469_ = pi087 & new_n409_ & pi132 & new_n442_;
  assign po41 = new_n552_ | new_n572_ | new_n520_ | new_n423_ | new_n469_;
  assign new_n471_ = pi087 & new_n409_ & pi133 & new_n442_;
  assign po42 = new_n553_ | new_n572_ | new_n521_ | new_n424_ | new_n471_;
  assign new_n473_ = pi087 & new_n409_ & pi134 & new_n442_;
  assign po43 = new_n554_ | new_n572_ | new_n522_ | new_n425_ | new_n473_;
  assign new_n475_ = pi087 & new_n409_ & pi135 & new_n442_;
  assign po44 = new_n555_ | new_n572_ | new_n523_ | new_n426_ | new_n475_;
  assign new_n477_ = pi087 & new_n409_ & pi136 & new_n442_;
  assign po45 = new_n556_ | new_n572_ | new_n524_ | new_n427_ | new_n477_;
  assign new_n479_ = pi087 & new_n409_ & pi137 & new_n442_;
  assign po46 = new_n557_ | new_n572_ | new_n525_ | new_n428_ | new_n479_;
  assign new_n481_ = pi087 & new_n409_ & pi138 & new_n442_;
  assign po47 = new_n558_ | new_n572_ | new_n526_ | new_n429_ | new_n481_;
  assign new_n483_ = pi087 & new_n409_ & pi139 & new_n442_;
  assign po48 = new_n559_ | new_n572_ | new_n527_ | new_n430_ | new_n483_;
  assign new_n485_ = pi087 & new_n409_ & pi140 & new_n442_;
  assign po49 = new_n560_ | new_n572_ | new_n528_ | new_n431_ | new_n485_;
  assign new_n487_ = pi087 & new_n409_ & pi141 & new_n442_;
  assign po50 = new_n561_ | new_n572_ | new_n529_ | new_n432_ | new_n487_;
  assign new_n489_ = pi087 & new_n409_ & pi142 & new_n442_;
  assign po51 = new_n562_ | new_n572_ | new_n530_ | new_n433_ | new_n489_;
  assign new_n491_ = pi087 & new_n409_ & pi143 & new_n442_;
  assign po52 = new_n563_ | new_n572_ | new_n531_ | new_n434_ | new_n491_;
  assign new_n493_ = pi087 & new_n409_ & pi144 & new_n442_;
  assign po53 = new_n564_ | new_n572_ | new_n532_ | new_n435_ | new_n493_;
  assign new_n495_ = pi087 & new_n409_ & pi145 & new_n442_;
  assign po54 = new_n565_ | new_n572_ | new_n533_ | new_n436_ | new_n495_;
  assign new_n497_ = pi087 & new_n409_ & pi146 & new_n442_;
  assign po55 = new_n566_ | new_n572_ | new_n534_ | new_n437_ | new_n497_;
  assign new_n499_ = pi087 & new_n409_ & pi147 & new_n442_;
  assign po56 = new_n567_ | new_n572_ | new_n535_ | new_n438_ | new_n499_;
  assign new_n501_ = pi087 & new_n409_ & pi148 & new_n442_;
  assign po57 = new_n568_ | new_n572_ | new_n536_ | new_n439_ | new_n501_;
  assign new_n503_ = pi087 & new_n409_ & pi149 & new_n442_;
  assign po58 = new_n569_ | new_n572_ | new_n537_ | new_n440_ | new_n503_;
  assign new_n505_ = pi087 & new_n409_ & pi150 & new_n442_;
  assign po59 = new_n570_ | new_n572_ | new_n538_ | new_n441_ | new_n505_;
  assign new_n507_ = pi087 & pi000 & pi151 & pi002;
  assign new_n508_ = pi087 & pi000 & pi152 & pi002;
  assign new_n509_ = pi087 & pi000 & pi153 & pi002;
  assign new_n510_ = pi087 & pi000 & pi154 & pi002;
  assign new_n511_ = pi087 & pi000 & pi155 & pi002;
  assign new_n512_ = pi087 & pi000 & pi156 & pi002;
  assign new_n513_ = pi087 & pi000 & pi157 & pi002;
  assign new_n514_ = pi087 & pi000 & pi158 & pi002;
  assign new_n515_ = pi087 & pi000 & pi159 & pi002;
  assign new_n516_ = pi087 & pi000 & pi160 & pi002;
  assign new_n517_ = pi087 & pi000 & pi161 & pi002;
  assign new_n518_ = pi087 & pi000 & pi162 & pi002;
  assign new_n519_ = pi087 & pi000 & pi163 & pi002;
  assign new_n520_ = pi087 & pi000 & pi164 & pi002;
  assign new_n521_ = pi087 & pi000 & pi165 & pi002;
  assign new_n522_ = pi087 & pi000 & pi166 & pi002;
  assign new_n523_ = pi087 & pi000 & pi167 & pi002;
  assign new_n524_ = pi087 & pi000 & pi168 & pi002;
  assign new_n525_ = pi087 & pi000 & pi169 & pi002;
  assign new_n526_ = pi087 & pi000 & pi170 & pi002;
  assign new_n527_ = pi087 & pi000 & pi171 & pi002;
  assign new_n528_ = pi087 & pi000 & pi172 & pi002;
  assign new_n529_ = pi087 & pi000 & pi173 & pi002;
  assign new_n530_ = pi087 & pi000 & pi174 & pi002;
  assign new_n531_ = pi087 & pi000 & pi175 & pi002;
  assign new_n532_ = pi087 & pi000 & pi176 & pi002;
  assign new_n533_ = pi087 & pi000 & pi177 & pi002;
  assign new_n534_ = pi087 & pi000 & pi178 & pi002;
  assign new_n535_ = pi087 & pi000 & pi179 & pi002;
  assign new_n536_ = pi087 & pi000 & pi180 & pi002;
  assign new_n537_ = pi087 & pi000 & pi181 & pi002;
  assign new_n538_ = pi087 & pi000 & pi182 & pi002;
  assign new_n539_ = pi087 & pi000 & new_n666_ & new_n442_;
  assign new_n540_ = pi087 & pi000 & new_n665_ & new_n442_;
  assign new_n541_ = pi087 & pi000 & new_n664_ & new_n442_;
  assign new_n542_ = pi087 & pi000 & new_n663_ & new_n442_;
  assign new_n543_ = pi087 & pi000 & new_n662_ & new_n442_;
  assign new_n544_ = pi087 & pi000 & new_n661_ & new_n442_;
  assign new_n545_ = pi087 & pi000 & new_n660_ & new_n442_;
  assign new_n546_ = pi087 & pi000 & new_n659_ & new_n442_;
  assign new_n547_ = pi087 & pi000 & new_n658_ & new_n442_;
  assign new_n548_ = pi087 & pi000 & new_n657_ & new_n442_;
  assign new_n549_ = pi087 & pi000 & new_n656_ & new_n442_;
  assign new_n550_ = pi087 & pi000 & new_n655_ & new_n442_;
  assign new_n551_ = pi087 & pi000 & new_n654_ & new_n442_;
  assign new_n552_ = pi087 & pi000 & new_n653_ & new_n442_;
  assign new_n553_ = pi087 & pi000 & new_n652_ & new_n442_;
  assign new_n554_ = pi087 & pi000 & new_n651_ & new_n442_;
  assign new_n555_ = pi087 & pi000 & new_n650_ & new_n442_;
  assign new_n556_ = pi087 & pi000 & new_n649_ & new_n442_;
  assign new_n557_ = pi087 & pi000 & new_n648_ & new_n442_;
  assign new_n558_ = pi087 & pi000 & new_n647_ & new_n442_;
  assign new_n559_ = pi087 & pi000 & new_n646_ & new_n442_;
  assign new_n560_ = pi087 & pi000 & new_n645_ & new_n442_;
  assign new_n561_ = pi087 & pi000 & new_n644_ & new_n442_;
  assign new_n562_ = pi087 & pi000 & new_n643_ & new_n442_;
  assign new_n563_ = pi087 & pi000 & new_n642_ & new_n442_;
  assign new_n564_ = pi087 & pi000 & new_n641_ & new_n442_;
  assign new_n565_ = pi087 & pi000 & new_n640_ & new_n442_;
  assign new_n566_ = pi087 & pi000 & new_n639_ & new_n442_;
  assign new_n567_ = pi087 & pi000 & new_n638_ & new_n442_;
  assign new_n568_ = pi087 & pi000 & new_n637_ & new_n442_;
  assign new_n569_ = pi087 & pi000 & new_n636_ & new_n442_;
  assign new_n570_ = pi087 & pi000 & new_n635_ & new_n442_;
  assign new_n571_ = ~pi087;
  assign new_n572_ = pi000 & new_n571_;
  assign new_n573_ = ~pi000;
  assign new_n574_ = pi184 & new_n573_ & pi183 & pi002;
  assign new_n575_ = pi184 & new_n573_ & pi185 & pi002;
  assign new_n576_ = pi184 & new_n573_ & pi186 & pi002;
  assign new_n577_ = pi184 & new_n573_ & pi187 & pi002;
  assign new_n578_ = ~pi002;
  assign new_n579_ = pi184 & new_n573_ & pi188 & new_n578_;
  assign po60 = new_n598_ | new_n579_;
  assign new_n581_ = pi184 & new_n573_ & pi189 & new_n578_;
  assign po61 = new_n593_ | new_n599_ | new_n606_ | new_n581_;
  assign new_n583_ = pi184 & new_n573_ & pi190 & new_n578_;
  assign po62 = new_n593_ | new_n600_ | new_n606_ | new_n583_;
  assign new_n585_ = pi184 & new_n573_ & pi191 & new_n578_;
  assign po63 = new_n601_ | new_n606_ | new_n594_ | new_n574_ | new_n585_;
  assign new_n587_ = pi184 & new_n573_ & pi192 & new_n578_;
  assign po64 = new_n602_ | new_n606_ | new_n595_ | new_n575_ | new_n587_;
  assign new_n589_ = pi184 & new_n573_ & pi193 & new_n578_;
  assign po65 = new_n603_ | new_n606_ | new_n596_ | new_n576_ | new_n589_;
  assign new_n591_ = pi184 & new_n573_ & pi194 & new_n578_;
  assign po66 = new_n604_ | new_n606_ | new_n597_ | new_n577_ | new_n591_;
  assign new_n593_ = pi002 & pi184 & pi000;
  assign new_n594_ = new_n593_ & pi195;
  assign new_n595_ = new_n593_ & pi196;
  assign new_n596_ = new_n593_ & pi197;
  assign new_n597_ = new_n593_ & pi198;
  assign new_n598_ = pi184 & pi000 & pi188 & new_n578_;
  assign new_n599_ = pi184 & pi000 & new_n672_ & new_n578_;
  assign new_n600_ = pi184 & pi000 & new_n671_ & new_n578_;
  assign new_n601_ = pi184 & pi000 & new_n670_ & new_n578_;
  assign new_n602_ = pi184 & pi000 & new_n669_ & new_n578_;
  assign new_n603_ = pi184 & pi000 & new_n668_ & new_n578_;
  assign new_n604_ = pi184 & pi000 & new_n667_ & new_n578_;
  assign new_n605_ = ~pi184;
  assign new_n606_ = pi000 & new_n605_;
  assign new_n607_ = ~pi057;
  assign new_n608_ = ~pi056;
  assign new_n609_ = ~pi055;
  assign new_n610_ = ~pi054;
  assign new_n611_ = ~pi053;
  assign new_n612_ = ~pi052;
  assign new_n613_ = ~pi051;
  assign new_n614_ = ~pi050;
  assign new_n615_ = ~pi049;
  assign new_n616_ = ~pi048;
  assign new_n617_ = ~pi047;
  assign new_n618_ = ~pi046;
  assign new_n619_ = ~pi045;
  assign new_n620_ = ~pi044;
  assign new_n621_ = ~pi043;
  assign new_n622_ = ~pi042;
  assign new_n623_ = ~pi041;
  assign new_n624_ = ~pi040;
  assign new_n625_ = ~pi039;
  assign new_n626_ = ~pi038;
  assign new_n627_ = ~pi037;
  assign new_n628_ = ~pi036;
  assign new_n629_ = ~pi035;
  assign new_n630_ = ~pi034;
  assign new_n631_ = ~pi033;
  assign new_n632_ = ~pi032;
  assign new_n633_ = ~pi031;
  assign new_n634_ = ~pi030;
  assign new_n635_ = ~pi150;
  assign new_n636_ = ~pi149;
  assign new_n637_ = ~pi148;
  assign new_n638_ = ~pi147;
  assign new_n639_ = ~pi146;
  assign new_n640_ = ~pi145;
  assign new_n641_ = ~pi144;
  assign new_n642_ = ~pi143;
  assign new_n643_ = ~pi142;
  assign new_n644_ = ~pi141;
  assign new_n645_ = ~pi140;
  assign new_n646_ = ~pi139;
  assign new_n647_ = ~pi138;
  assign new_n648_ = ~pi137;
  assign new_n649_ = ~pi136;
  assign new_n650_ = ~pi135;
  assign new_n651_ = ~pi134;
  assign new_n652_ = ~pi133;
  assign new_n653_ = ~pi132;
  assign new_n654_ = ~pi131;
  assign new_n655_ = ~pi130;
  assign new_n656_ = ~pi129;
  assign new_n657_ = ~pi128;
  assign new_n658_ = ~pi127;
  assign new_n659_ = ~pi126;
  assign new_n660_ = ~pi125;
  assign new_n661_ = ~pi124;
  assign new_n662_ = ~pi123;
  assign new_n663_ = ~pi122;
  assign new_n664_ = ~pi121;
  assign new_n665_ = ~pi120;
  assign new_n666_ = ~pi119;
  assign new_n667_ = ~pi194;
  assign new_n668_ = ~pi193;
  assign new_n669_ = ~pi192;
  assign new_n670_ = ~pi191;
  assign new_n671_ = ~pi190;
  assign new_n672_ = ~pi189;
endmodule


