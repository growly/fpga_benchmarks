// Benchmark "i6" written by ABC on Thu Mar 19 13:02:36 2020

module i6 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47,
    po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46,
    po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58,
    po59, po60, po61, po62, po63, po64, po65, po66;
  wire new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_,
    new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n238_, new_n240_, new_n242_, new_n244_, new_n246_,
    new_n248_, new_n250_, new_n252_, new_n254_, new_n256_, new_n258_,
    new_n260_, new_n262_, new_n264_, new_n266_, new_n268_, new_n270_,
    new_n272_, new_n274_, new_n276_, new_n278_, new_n280_, new_n282_,
    new_n284_, new_n286_, new_n288_, new_n290_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n356_, new_n358_, new_n360_, new_n362_, new_n364_,
    new_n366_, new_n368_, new_n370_, new_n372_, new_n374_, new_n376_,
    new_n378_, new_n380_, new_n382_, new_n384_, new_n386_, new_n388_,
    new_n390_, new_n392_, new_n394_, new_n396_, new_n398_, new_n400_,
    new_n402_, new_n404_, new_n406_, new_n408_, new_n410_, new_n412_,
    new_n414_, new_n416_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n463_, new_n465_,
    new_n467_, new_n469_, new_n471_, new_n473_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_;
  assign new_n206_ = ~pi000;
  assign new_n207_ = ~pi001;
  assign new_n208_ = new_n206_ & pi002 & new_n207_;
  assign new_n209_ = new_n206_ & pi003 & new_n207_;
  assign new_n210_ = new_n206_ & pi004 & new_n207_;
  assign new_n211_ = new_n206_ & pi005 & new_n207_;
  assign new_n212_ = new_n206_ & pi006 & new_n207_;
  assign new_n213_ = new_n206_ & pi007 & new_n207_;
  assign new_n214_ = new_n206_ & pi008 & new_n207_;
  assign new_n215_ = new_n206_ & pi009 & new_n207_;
  assign new_n216_ = new_n206_ & pi010 & new_n207_;
  assign new_n217_ = new_n206_ & pi011 & new_n207_;
  assign new_n218_ = new_n206_ & pi012 & new_n207_;
  assign new_n219_ = new_n206_ & pi013 & new_n207_;
  assign new_n220_ = new_n206_ & pi014 & new_n207_;
  assign new_n221_ = new_n206_ & pi015 & new_n207_;
  assign new_n222_ = new_n206_ & pi016 & new_n207_;
  assign new_n223_ = new_n206_ & pi017 & new_n207_;
  assign new_n224_ = new_n206_ & pi018 & new_n207_;
  assign new_n225_ = new_n206_ & pi019 & new_n207_;
  assign new_n226_ = new_n206_ & pi020 & new_n207_;
  assign new_n227_ = new_n206_ & pi021 & new_n207_;
  assign new_n228_ = new_n206_ & pi022 & new_n207_;
  assign new_n229_ = new_n206_ & pi023 & new_n207_;
  assign new_n230_ = new_n206_ & pi024 & new_n207_;
  assign new_n231_ = new_n206_ & pi025 & new_n207_;
  assign new_n232_ = new_n206_ & pi026 & new_n207_;
  assign new_n233_ = new_n206_ & pi027 & new_n207_;
  assign new_n234_ = new_n206_ & pi028 & new_n207_;
  assign new_n235_ = new_n206_ & pi029 & new_n207_;
  assign new_n236_ = pi000 & pi030 & new_n207_;
  assign po00 = new_n292_ | new_n208_ | new_n236_;
  assign new_n238_ = pi000 & pi031 & new_n207_;
  assign po01 = new_n293_ | new_n209_ | new_n238_;
  assign new_n240_ = pi000 & pi032 & new_n207_;
  assign po02 = new_n294_ | new_n210_ | new_n240_;
  assign new_n242_ = pi000 & pi033 & new_n207_;
  assign po03 = new_n295_ | new_n211_ | new_n242_;
  assign new_n244_ = pi000 & pi034 & new_n207_;
  assign po04 = new_n296_ | new_n212_ | new_n244_;
  assign new_n246_ = pi000 & pi035 & new_n207_;
  assign po05 = new_n297_ | new_n213_ | new_n246_;
  assign new_n248_ = pi000 & pi036 & new_n207_;
  assign po06 = new_n298_ | new_n214_ | new_n248_;
  assign new_n250_ = pi000 & pi037 & new_n207_;
  assign po07 = new_n299_ | new_n215_ | new_n250_;
  assign new_n252_ = pi000 & pi038 & new_n207_;
  assign po08 = new_n300_ | new_n216_ | new_n252_;
  assign new_n254_ = pi000 & pi039 & new_n207_;
  assign po09 = new_n301_ | new_n217_ | new_n254_;
  assign new_n256_ = pi000 & pi040 & new_n207_;
  assign po10 = new_n302_ | new_n218_ | new_n256_;
  assign new_n258_ = pi000 & pi041 & new_n207_;
  assign po11 = new_n303_ | new_n219_ | new_n258_;
  assign new_n260_ = pi000 & pi042 & new_n207_;
  assign po12 = new_n304_ | new_n220_ | new_n260_;
  assign new_n262_ = pi000 & pi043 & new_n207_;
  assign po13 = new_n305_ | new_n221_ | new_n262_;
  assign new_n264_ = pi000 & pi044 & new_n207_;
  assign po14 = new_n306_ | new_n222_ | new_n264_;
  assign new_n266_ = pi000 & pi045 & new_n207_;
  assign po15 = new_n307_ | new_n223_ | new_n266_;
  assign new_n268_ = pi000 & pi046 & new_n207_;
  assign po16 = new_n308_ | new_n224_ | new_n268_;
  assign new_n270_ = pi000 & pi047 & new_n207_;
  assign po17 = new_n309_ | new_n225_ | new_n270_;
  assign new_n272_ = pi000 & pi048 & new_n207_;
  assign po18 = new_n310_ | new_n226_ | new_n272_;
  assign new_n274_ = pi000 & pi049 & new_n207_;
  assign po19 = new_n311_ | new_n227_ | new_n274_;
  assign new_n276_ = pi000 & pi050 & new_n207_;
  assign po20 = new_n312_ | new_n228_ | new_n276_;
  assign new_n278_ = pi000 & pi051 & new_n207_;
  assign po21 = new_n313_ | new_n229_ | new_n278_;
  assign new_n280_ = pi000 & pi052 & new_n207_;
  assign po22 = new_n314_ | new_n230_ | new_n280_;
  assign new_n282_ = pi000 & pi053 & new_n207_;
  assign po23 = new_n315_ | new_n231_ | new_n282_;
  assign new_n284_ = pi000 & pi054 & new_n207_;
  assign po24 = new_n316_ | new_n232_ | new_n284_;
  assign new_n286_ = pi000 & pi055 & new_n207_;
  assign po25 = new_n317_ | new_n233_ | new_n286_;
  assign new_n288_ = pi000 & pi056 & new_n207_;
  assign po26 = new_n318_ | new_n234_ | new_n288_;
  assign new_n290_ = pi000 & pi057 & new_n207_;
  assign po27 = new_n319_ | new_n235_ | new_n290_;
  assign new_n292_ = pi000 & new_n511_ & pi001;
  assign new_n293_ = pi000 & new_n510_ & pi001;
  assign new_n294_ = pi000 & new_n509_ & pi001;
  assign new_n295_ = pi000 & new_n508_ & pi001;
  assign new_n296_ = pi000 & new_n507_ & pi001;
  assign new_n297_ = pi000 & new_n506_ & pi001;
  assign new_n298_ = pi000 & new_n505_ & pi001;
  assign new_n299_ = pi000 & new_n504_ & pi001;
  assign new_n300_ = pi000 & new_n503_ & pi001;
  assign new_n301_ = pi000 & new_n502_ & pi001;
  assign new_n302_ = pi000 & new_n501_ & pi001;
  assign new_n303_ = pi000 & new_n500_ & pi001;
  assign new_n304_ = pi000 & new_n499_ & pi001;
  assign new_n305_ = pi000 & new_n498_ & pi001;
  assign new_n306_ = pi000 & new_n497_ & pi001;
  assign new_n307_ = pi000 & new_n496_ & pi001;
  assign new_n308_ = pi000 & new_n495_ & pi001;
  assign new_n309_ = pi000 & new_n494_ & pi001;
  assign new_n310_ = pi000 & new_n493_ & pi001;
  assign new_n311_ = pi000 & new_n492_ & pi001;
  assign new_n312_ = pi000 & new_n491_ & pi001;
  assign new_n313_ = pi000 & new_n490_ & pi001;
  assign new_n314_ = pi000 & new_n489_ & pi001;
  assign new_n315_ = pi000 & new_n488_ & pi001;
  assign new_n316_ = pi000 & new_n487_ & pi001;
  assign new_n317_ = pi000 & new_n486_ & pi001;
  assign new_n318_ = pi000 & new_n485_ & pi001;
  assign new_n319_ = pi000 & new_n484_ & pi001;
  assign new_n320_ = ~pi000;
  assign new_n321_ = ~pi001;
  assign new_n322_ = pi059 & new_n321_ & pi058 & new_n320_;
  assign new_n323_ = pi059 & new_n321_ & pi060 & new_n320_;
  assign new_n324_ = pi059 & new_n321_ & pi061 & new_n320_;
  assign new_n325_ = pi059 & new_n321_ & pi062 & new_n320_;
  assign new_n326_ = pi059 & new_n321_ & pi063 & new_n320_;
  assign new_n327_ = pi059 & new_n321_ & pi064 & new_n320_;
  assign new_n328_ = pi059 & new_n321_ & pi065 & new_n320_;
  assign new_n329_ = pi059 & new_n321_ & pi066 & new_n320_;
  assign new_n330_ = pi059 & new_n321_ & pi067 & new_n320_;
  assign new_n331_ = pi059 & new_n321_ & pi068 & new_n320_;
  assign new_n332_ = pi059 & new_n321_ & pi069 & new_n320_;
  assign new_n333_ = pi059 & new_n321_ & pi070 & new_n320_;
  assign new_n334_ = pi059 & new_n321_ & pi071 & new_n320_;
  assign new_n335_ = pi059 & new_n321_ & pi072 & new_n320_;
  assign new_n336_ = pi059 & new_n321_ & pi073 & new_n320_;
  assign new_n337_ = pi059 & new_n321_ & pi074 & new_n320_;
  assign new_n338_ = pi059 & new_n321_ & pi075 & new_n320_;
  assign new_n339_ = pi059 & new_n321_ & pi076 & new_n320_;
  assign new_n340_ = pi059 & new_n321_ & pi077 & new_n320_;
  assign new_n341_ = pi059 & new_n321_ & pi078 & new_n320_;
  assign new_n342_ = pi059 & new_n321_ & pi079 & new_n320_;
  assign new_n343_ = pi059 & new_n321_ & pi080 & new_n320_;
  assign new_n344_ = pi059 & new_n321_ & pi081 & new_n320_;
  assign new_n345_ = pi059 & new_n321_ & pi082 & new_n320_;
  assign new_n346_ = pi059 & new_n321_ & pi083 & new_n320_;
  assign new_n347_ = pi059 & new_n321_ & pi084 & new_n320_;
  assign new_n348_ = pi059 & new_n321_ & pi085 & new_n320_;
  assign new_n349_ = pi059 & new_n321_ & pi086 & new_n320_;
  assign new_n350_ = pi059 & new_n321_ & pi087 & new_n320_;
  assign new_n351_ = pi059 & new_n321_ & pi088 & new_n320_;
  assign new_n352_ = pi059 & new_n321_ & pi089 & new_n320_;
  assign new_n353_ = pi059 & new_n321_ & pi090 & new_n320_;
  assign new_n354_ = pi059 & new_n321_ & pi091 & pi000;
  assign po28 = new_n322_ | new_n354_ | new_n418_ | new_n451_;
  assign new_n356_ = pi059 & new_n321_ & pi092 & pi000;
  assign po29 = new_n323_ | new_n356_ | new_n419_ | new_n451_;
  assign new_n358_ = pi059 & new_n321_ & pi093 & pi000;
  assign po30 = new_n324_ | new_n358_ | new_n420_ | new_n451_;
  assign new_n360_ = pi059 & new_n321_ & pi094 & pi000;
  assign po31 = new_n325_ | new_n360_ | new_n421_ | new_n451_;
  assign new_n362_ = pi059 & new_n321_ & pi095 & pi000;
  assign po32 = new_n326_ | new_n362_ | new_n422_ | new_n451_;
  assign new_n364_ = pi059 & new_n321_ & pi096 & pi000;
  assign po33 = new_n327_ | new_n364_ | new_n423_ | new_n451_;
  assign new_n366_ = pi059 & new_n321_ & pi097 & pi000;
  assign po34 = new_n328_ | new_n366_ | new_n424_ | new_n451_;
  assign new_n368_ = pi059 & new_n321_ & pi098 & pi000;
  assign po35 = new_n329_ | new_n368_ | new_n425_ | new_n451_;
  assign new_n370_ = pi059 & new_n321_ & pi099 & pi000;
  assign po36 = new_n330_ | new_n370_ | new_n426_ | new_n451_;
  assign new_n372_ = pi059 & new_n321_ & pi100 & pi000;
  assign po37 = new_n331_ | new_n372_ | new_n427_ | new_n451_;
  assign new_n374_ = pi059 & new_n321_ & pi101 & pi000;
  assign po38 = new_n332_ | new_n374_ | new_n428_ | new_n451_;
  assign new_n376_ = pi059 & new_n321_ & pi102 & pi000;
  assign po39 = new_n333_ | new_n376_ | new_n429_ | new_n451_;
  assign new_n378_ = pi059 & new_n321_ & pi103 & pi000;
  assign po40 = new_n334_ | new_n378_ | new_n430_ | new_n451_;
  assign new_n380_ = pi059 & new_n321_ & pi104 & pi000;
  assign po41 = new_n335_ | new_n380_ | new_n431_ | new_n451_;
  assign new_n382_ = pi059 & new_n321_ & pi105 & pi000;
  assign po42 = new_n336_ | new_n382_ | new_n432_ | new_n451_;
  assign new_n384_ = pi059 & new_n321_ & pi106 & pi000;
  assign po43 = new_n337_ | new_n384_ | new_n433_ | new_n451_;
  assign new_n386_ = pi059 & new_n321_ & pi107 & pi000;
  assign po44 = new_n338_ | new_n386_ | new_n434_ | new_n451_;
  assign new_n388_ = pi059 & new_n321_ & pi108 & pi000;
  assign po45 = new_n339_ | new_n388_ | new_n435_ | new_n451_;
  assign new_n390_ = pi059 & new_n321_ & pi109 & pi000;
  assign po46 = new_n340_ | new_n390_ | new_n436_ | new_n451_;
  assign new_n392_ = pi059 & new_n321_ & pi110 & pi000;
  assign po47 = new_n341_ | new_n392_ | new_n437_ | new_n451_;
  assign new_n394_ = pi059 & new_n321_ & pi111 & pi000;
  assign po48 = new_n342_ | new_n394_ | new_n438_ | new_n451_;
  assign new_n396_ = pi059 & new_n321_ & pi112 & pi000;
  assign po49 = new_n343_ | new_n396_ | new_n439_ | new_n451_;
  assign new_n398_ = pi059 & new_n321_ & pi113 & pi000;
  assign po50 = new_n344_ | new_n398_ | new_n440_ | new_n451_;
  assign new_n400_ = pi059 & new_n321_ & pi114 & pi000;
  assign po51 = new_n345_ | new_n400_ | new_n441_ | new_n451_;
  assign new_n402_ = pi059 & new_n321_ & pi115 & pi000;
  assign po52 = new_n346_ | new_n402_ | new_n442_ | new_n451_;
  assign new_n404_ = pi059 & new_n321_ & pi116 & pi000;
  assign po53 = new_n347_ | new_n404_ | new_n443_ | new_n451_;
  assign new_n406_ = pi059 & new_n321_ & pi117 & pi000;
  assign po54 = new_n348_ | new_n406_ | new_n444_ | new_n451_;
  assign new_n408_ = pi059 & new_n321_ & pi118 & pi000;
  assign po55 = new_n349_ | new_n408_ | new_n445_ | new_n451_;
  assign new_n410_ = pi059 & new_n321_ & pi119 & pi000;
  assign po56 = new_n350_ | new_n410_ | new_n446_ | new_n451_;
  assign new_n412_ = pi059 & new_n321_ & pi120 & pi000;
  assign po57 = new_n351_ | new_n412_ | new_n447_ | new_n451_;
  assign new_n414_ = pi059 & new_n321_ & pi121 & pi000;
  assign po58 = new_n352_ | new_n414_ | new_n448_ | new_n451_;
  assign new_n416_ = pi059 & new_n321_ & pi122 & pi000;
  assign po59 = new_n353_ | new_n416_ | new_n449_ | new_n451_;
  assign new_n418_ = pi059 & pi001 & new_n543_ & pi000;
  assign new_n419_ = pi059 & pi001 & new_n542_ & pi000;
  assign new_n420_ = pi059 & pi001 & new_n541_ & pi000;
  assign new_n421_ = pi059 & pi001 & new_n540_ & pi000;
  assign new_n422_ = pi059 & pi001 & new_n539_ & pi000;
  assign new_n423_ = pi059 & pi001 & new_n538_ & pi000;
  assign new_n424_ = pi059 & pi001 & new_n537_ & pi000;
  assign new_n425_ = pi059 & pi001 & new_n536_ & pi000;
  assign new_n426_ = pi059 & pi001 & new_n535_ & pi000;
  assign new_n427_ = pi059 & pi001 & new_n534_ & pi000;
  assign new_n428_ = pi059 & pi001 & new_n533_ & pi000;
  assign new_n429_ = pi059 & pi001 & new_n532_ & pi000;
  assign new_n430_ = pi059 & pi001 & new_n531_ & pi000;
  assign new_n431_ = pi059 & pi001 & new_n530_ & pi000;
  assign new_n432_ = pi059 & pi001 & new_n529_ & pi000;
  assign new_n433_ = pi059 & pi001 & new_n528_ & pi000;
  assign new_n434_ = pi059 & pi001 & new_n527_ & pi000;
  assign new_n435_ = pi059 & pi001 & new_n526_ & pi000;
  assign new_n436_ = pi059 & pi001 & new_n525_ & pi000;
  assign new_n437_ = pi059 & pi001 & new_n524_ & pi000;
  assign new_n438_ = pi059 & pi001 & new_n523_ & pi000;
  assign new_n439_ = pi059 & pi001 & new_n522_ & pi000;
  assign new_n440_ = pi059 & pi001 & new_n521_ & pi000;
  assign new_n441_ = pi059 & pi001 & new_n520_ & pi000;
  assign new_n442_ = pi059 & pi001 & new_n519_ & pi000;
  assign new_n443_ = pi059 & pi001 & new_n518_ & pi000;
  assign new_n444_ = pi059 & pi001 & new_n517_ & pi000;
  assign new_n445_ = pi059 & pi001 & new_n516_ & pi000;
  assign new_n446_ = pi059 & pi001 & new_n515_ & pi000;
  assign new_n447_ = pi059 & pi001 & new_n514_ & pi000;
  assign new_n448_ = pi059 & pi001 & new_n513_ & pi000;
  assign new_n449_ = pi059 & pi001 & new_n512_ & pi000;
  assign new_n450_ = ~pi059;
  assign new_n451_ = pi001 & new_n450_;
  assign new_n452_ = ~pi000;
  assign new_n453_ = ~pi001;
  assign new_n454_ = pi124 & new_n453_ & pi123 & new_n452_;
  assign new_n455_ = pi124 & new_n453_ & pi125 & new_n452_;
  assign new_n456_ = pi124 & new_n453_ & pi126 & new_n452_;
  assign new_n457_ = pi124 & new_n453_ & pi127 & new_n452_;
  assign new_n458_ = pi124 & new_n453_ & pi128 & new_n452_;
  assign new_n459_ = pi124 & new_n453_ & pi129 & new_n452_;
  assign new_n460_ = pi124 & new_n453_ & pi130 & new_n452_;
  assign new_n461_ = pi124 & new_n453_ & pi131 & pi000;
  assign po60 = new_n475_ | new_n454_ | new_n461_;
  assign new_n463_ = pi124 & new_n453_ & pi132 & pi000;
  assign po61 = new_n455_ | new_n463_ | new_n476_ | new_n483_;
  assign new_n465_ = pi124 & new_n453_ & pi133 & pi000;
  assign po62 = new_n456_ | new_n465_ | new_n477_ | new_n483_;
  assign new_n467_ = pi124 & new_n453_ & pi134 & pi000;
  assign po63 = new_n457_ | new_n467_ | new_n478_ | new_n483_;
  assign new_n469_ = pi124 & new_n453_ & pi135 & pi000;
  assign po64 = new_n458_ | new_n469_ | new_n479_ | new_n483_;
  assign new_n471_ = pi124 & new_n453_ & pi136 & pi000;
  assign po65 = new_n459_ | new_n471_ | new_n480_ | new_n483_;
  assign new_n473_ = pi124 & new_n453_ & pi137 & pi000;
  assign po66 = new_n460_ | new_n473_ | new_n481_ | new_n483_;
  assign new_n475_ = pi124 & pi001 & pi131 & pi000;
  assign new_n476_ = pi124 & pi001 & new_n549_ & pi000;
  assign new_n477_ = pi124 & pi001 & new_n548_ & pi000;
  assign new_n478_ = pi124 & pi001 & new_n547_ & pi000;
  assign new_n479_ = pi124 & pi001 & new_n546_ & pi000;
  assign new_n480_ = pi124 & pi001 & new_n545_ & pi000;
  assign new_n481_ = pi124 & pi001 & new_n544_ & pi000;
  assign new_n482_ = ~pi124;
  assign new_n483_ = pi001 & new_n482_;
  assign new_n484_ = ~pi057;
  assign new_n485_ = ~pi056;
  assign new_n486_ = ~pi055;
  assign new_n487_ = ~pi054;
  assign new_n488_ = ~pi053;
  assign new_n489_ = ~pi052;
  assign new_n490_ = ~pi051;
  assign new_n491_ = ~pi050;
  assign new_n492_ = ~pi049;
  assign new_n493_ = ~pi048;
  assign new_n494_ = ~pi047;
  assign new_n495_ = ~pi046;
  assign new_n496_ = ~pi045;
  assign new_n497_ = ~pi044;
  assign new_n498_ = ~pi043;
  assign new_n499_ = ~pi042;
  assign new_n500_ = ~pi041;
  assign new_n501_ = ~pi040;
  assign new_n502_ = ~pi039;
  assign new_n503_ = ~pi038;
  assign new_n504_ = ~pi037;
  assign new_n505_ = ~pi036;
  assign new_n506_ = ~pi035;
  assign new_n507_ = ~pi034;
  assign new_n508_ = ~pi033;
  assign new_n509_ = ~pi032;
  assign new_n510_ = ~pi031;
  assign new_n511_ = ~pi030;
  assign new_n512_ = ~pi122;
  assign new_n513_ = ~pi121;
  assign new_n514_ = ~pi120;
  assign new_n515_ = ~pi119;
  assign new_n516_ = ~pi118;
  assign new_n517_ = ~pi117;
  assign new_n518_ = ~pi116;
  assign new_n519_ = ~pi115;
  assign new_n520_ = ~pi114;
  assign new_n521_ = ~pi113;
  assign new_n522_ = ~pi112;
  assign new_n523_ = ~pi111;
  assign new_n524_ = ~pi110;
  assign new_n525_ = ~pi109;
  assign new_n526_ = ~pi108;
  assign new_n527_ = ~pi107;
  assign new_n528_ = ~pi106;
  assign new_n529_ = ~pi105;
  assign new_n530_ = ~pi104;
  assign new_n531_ = ~pi103;
  assign new_n532_ = ~pi102;
  assign new_n533_ = ~pi101;
  assign new_n534_ = ~pi100;
  assign new_n535_ = ~pi099;
  assign new_n536_ = ~pi098;
  assign new_n537_ = ~pi097;
  assign new_n538_ = ~pi096;
  assign new_n539_ = ~pi095;
  assign new_n540_ = ~pi094;
  assign new_n541_ = ~pi093;
  assign new_n542_ = ~pi092;
  assign new_n543_ = ~pi091;
  assign new_n544_ = ~pi137;
  assign new_n545_ = ~pi136;
  assign new_n546_ = ~pi135;
  assign new_n547_ = ~pi134;
  assign new_n548_ = ~pi133;
  assign new_n549_ = ~pi132;
endmodule


