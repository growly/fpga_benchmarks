// Benchmark "i10" written by ABC on Thu Mar 19 13:02:36 2020

module i10 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255, pi256,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223;
  wire new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n532_, new_n534_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n591_, new_n592_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n652_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n697_, new_n699_,
    new_n701_, new_n703_, new_n705_, new_n707_, new_n709_, new_n711_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n918_, new_n919_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1052_, new_n1053_, new_n1054_,
    new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_,
    new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_,
    new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_,
    new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_,
    new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_,
    new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_,
    new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_,
    new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_,
    new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_,
    new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_,
    new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_,
    new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_,
    new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_,
    new_n1272_, new_n1273_, new_n1274_, new_n1276_, new_n1278_, new_n1280_,
    new_n1282_, new_n1284_, new_n1286_, new_n1288_, new_n1290_, new_n1292_,
    new_n1294_, new_n1296_, new_n1298_, new_n1299_, new_n1300_, new_n1301_,
    new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_,
    new_n1308_, new_n1310_, new_n1312_, new_n1314_, new_n1316_, new_n1318_,
    new_n1320_, new_n1322_, new_n1324_, new_n1326_, new_n1328_, new_n1329_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_,
    new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1352_, new_n1353_,
    new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1359_, new_n1360_,
    new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1366_, new_n1367_,
    new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1374_,
    new_n1376_, new_n1378_, new_n1380_, new_n1382_, new_n1383_, new_n1384_,
    new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_,
    new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_,
    new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_,
    new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_,
    new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_,
    new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_,
    new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_,
    new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_,
    new_n1433_, new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1440_,
    new_n1441_, new_n1443_, new_n1445_, new_n1447_, new_n1449_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1457_, new_n1458_, new_n1459_,
    new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_,
    new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_,
    new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_,
    new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1488_, new_n1489_, new_n1491_,
    new_n1494_, new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_,
    new_n1502_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1516_,
    new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_,
    new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_,
    new_n1530_, new_n1532_, new_n1533_, new_n1535_, new_n1536_, new_n1537_,
    new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_,
    new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_,
    new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1557_, new_n1558_,
    new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_,
    new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_,
    new_n1573_, new_n1575_, new_n1577_, new_n1578_, new_n1579_, new_n1580_,
    new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_,
    new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_,
    new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_,
    new_n1599_, new_n1602_, new_n1604_, new_n1605_, new_n1606_, new_n1607_,
    new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_,
    new_n1615_, new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_,
    new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_,
    new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_,
    new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_,
    new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_,
    new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_,
    new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_,
    new_n1661_, new_n1662_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_,
    new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1680_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1687_,
    new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_,
    new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_,
    new_n1700_, new_n1701_, new_n1702_, new_n1704_, new_n1706_, new_n1707_,
    new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1714_,
    new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_,
    new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_,
    new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_,
    new_n1734_, new_n1736_, new_n1738_, new_n1740_, new_n1742_, new_n1744_,
    new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_,
    new_n1752_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1765_,
    new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1771_, new_n1772_,
    new_n1773_, new_n1774_, new_n1776_, new_n1777_, new_n1778_, new_n1780_,
    new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_,
    new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1795_, new_n1796_,
    new_n1797_, new_n1798_, new_n1800_, new_n1802_, new_n1803_, new_n1804_,
    new_n1806_, new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1821_, new_n1823_, new_n1825_, new_n1827_, new_n1829_,
    new_n1831_, new_n1833_, new_n1835_, new_n1837_, new_n1839_, new_n1840_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1874_,
    new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_,
    new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_,
    new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_,
    new_n1893_, new_n1894_, new_n1895_, new_n1902_, new_n1903_, new_n1904_,
    new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1911_,
    new_n1913_, new_n1915_, new_n1917_, new_n1919_, new_n1921_, new_n1922_,
    new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_,
    new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_,
    new_n1935_, new_n1936_, new_n1937_, new_n1939_, new_n1940_, new_n1942_,
    new_n1944_, new_n1946_, new_n1948_, new_n1950_, new_n1953_, new_n1954_,
    new_n1955_, new_n1956_, new_n1958_, new_n1960_, new_n1961_, new_n1962_,
    new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1968_, new_n1969_,
    new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_,
    new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_,
    new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1988_,
    new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_,
    new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_,
    new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_,
    new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_,
    new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_,
    new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_,
    new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_,
    new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_,
    new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_,
    new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_,
    new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_,
    new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_,
    new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_,
    new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_,
    new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_,
    new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_,
    new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2091_,
    new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_,
    new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_,
    new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_,
    new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_,
    new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_,
    new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_,
    new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_,
    new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_,
    new_n2140_, new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_,
    new_n2146_, new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2151_,
    new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_,
    new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_,
    new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_,
    new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_,
    new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_,
    new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_,
    new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_,
    new_n2194_, new_n2195_, new_n2196_, new_n2197_, new_n2198_, new_n2199_,
    new_n2200_, new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2205_,
    new_n2206_, new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_,
    new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2217_,
    new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_, new_n2223_,
    new_n2224_, new_n2225_, new_n2226_, new_n2227_, new_n2228_, new_n2229_,
    new_n2230_, new_n2231_, new_n2232_, new_n2233_, new_n2234_, new_n2235_,
    new_n2236_, new_n2237_, new_n2238_, new_n2239_, new_n2240_, new_n2241_,
    new_n2242_, new_n2243_, new_n2244_, new_n2245_, new_n2246_, new_n2247_,
    new_n2248_, new_n2249_, new_n2250_, new_n2251_, new_n2252_, new_n2253_,
    new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2258_, new_n2259_,
    new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_, new_n2265_,
    new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_, new_n2271_,
    new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_, new_n2277_,
    new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_, new_n2283_,
    new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_, new_n2289_,
    new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_, new_n2295_,
    new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_, new_n2301_,
    new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_, new_n2307_,
    new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_, new_n2313_,
    new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_, new_n2319_,
    new_n2320_, new_n2321_, new_n2322_, new_n2324_, new_n2325_, new_n2326_,
    new_n2327_, new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2334_,
    new_n2335_, new_n2336_, new_n2337_, new_n2339_, new_n2340_, new_n2341_,
    new_n2342_, new_n2344_, new_n2345_, new_n2346_, new_n2347_, new_n2349_,
    new_n2350_, new_n2351_, new_n2352_, new_n2354_, new_n2355_, new_n2356_,
    new_n2357_, new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_,
    new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_,
    new_n2369_, new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_,
    new_n2375_, new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_,
    new_n2381_, new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_,
    new_n2387_, new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_,
    new_n2393_, new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_,
    new_n2399_, new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_,
    new_n2405_, new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_,
    new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_,
    new_n2417_, new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_,
    new_n2423_, new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_,
    new_n2429_, new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_,
    new_n2435_, new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_,
    new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_,
    new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_,
    new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_,
    new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_,
    new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_,
    new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_,
    new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_,
    new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_,
    new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_,
    new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_,
    new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_,
    new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_,
    new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_,
    new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_,
    new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_,
    new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_,
    new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_,
    new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_,
    new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_,
    new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_,
    new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_,
    new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_,
    new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_,
    new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_,
    new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_,
    new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_,
    new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_,
    new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_,
    new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_,
    new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_,
    new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_,
    new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_,
    new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_,
    new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_,
    new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_,
    new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_,
    new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_,
    new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_,
    new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2674_, new_n2675_,
    new_n2676_, new_n2677_, new_n2679_, new_n2680_, new_n2681_, new_n2682_,
    new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2689_, new_n2690_,
    new_n2691_, new_n2692_, new_n2694_, new_n2695_, new_n2696_, new_n2697_,
    new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_,
    new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_,
    new_n2710_, new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_,
    new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_,
    new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_,
    new_n2728_, new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_,
    new_n2734_, new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_,
    new_n2740_, new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_,
    new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_,
    new_n2752_, new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_,
    new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_,
    new_n2764_, new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2769_,
    new_n2770_, new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_,
    new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_,
    new_n2782_, new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_,
    new_n2788_, new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_,
    new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_,
    new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_,
    new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_,
    new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_,
    new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_,
    new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_,
    new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_,
    new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_,
    new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_,
    new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_,
    new_n2854_, new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_,
    new_n2860_, new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_,
    new_n2866_, new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_,
    new_n2872_, new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_,
    new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_,
    new_n2884_, new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_,
    new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_,
    new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_,
    new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_,
    new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_,
    new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_,
    new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_,
    new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_,
    new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_,
    new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_,
    new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_, new_n2949_,
    new_n2950_, new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_,
    new_n2956_, new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_,
    new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_,
    new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_,
    new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_;
  assign po000 = ~po091;
  assign new_n483_ = ~new_n2258_;
  assign new_n484_ = new_n483_ & pi000;
  assign new_n485_ = ~new_n2253_;
  assign new_n486_ = ~new_n2218_;
  assign new_n487_ = new_n485_ & new_n486_ & pi001;
  assign new_n488_ = ~new_n2248_;
  assign new_n489_ = ~new_n2223_;
  assign new_n490_ = new_n486_ & pi002 & new_n489_ & new_n488_;
  assign new_n491_ = ~new_n2233_;
  assign new_n492_ = ~new_n2228_;
  assign new_n493_ = new_n489_ & new_n491_ & pi003 & new_n492_ & new_n486_;
  assign new_n494_ = new_n484_ | new_n490_ | new_n493_ | new_n487_;
  assign new_n495_ = ~new_n1540_;
  assign new_n496_ = ~new_n828_;
  assign new_n497_ = new_n495_ & new_n877_ & new_n496_ & pi004;
  assign new_n498_ = po065 & new_n854_;
  assign new_n499_ = new_n2007_ & po065;
  assign new_n500_ = ~new_n497_;
  assign new_n501_ = ~po065;
  assign new_n502_ = ~pi005;
  assign new_n503_ = pi004 & new_n892_;
  assign new_n504_ = ~new_n503_;
  assign new_n505_ = new_n592_ & new_n1719_;
  assign new_n506_ = new_n1032_ & new_n1719_ & new_n1026_;
  assign new_n507_ = new_n1020_ & new_n1719_ & new_n1014_;
  assign new_n508_ = new_n1008_ & new_n1719_ & new_n1002_;
  assign new_n509_ = new_n996_ & new_n1719_ & new_n990_;
  assign new_n510_ = new_n984_ & new_n1719_ & new_n978_;
  assign new_n511_ = new_n972_ & new_n1719_ & new_n966_;
  assign new_n512_ = new_n1044_ & new_n1719_ & new_n1043_;
  assign new_n513_ = new_n1042_ & new_n1719_ & new_n1041_;
  assign po001 = new_n1026_ & new_n1002_ & new_n978_ & new_n1043_ & new_n1041_ & new_n966_ & new_n990_ & new_n505_ & new_n1014_;
  assign po002 = new_n1032_ & new_n1008_ & new_n984_ & new_n1044_ & new_n1042_ & new_n972_ & new_n996_ & new_n1719_ & new_n1020_;
  assign new_n516_ = new_n1026_ & new_n1014_ & new_n1002_ & new_n990_ & new_n996_ & new_n1008_ & new_n1032_ & new_n1020_;
  assign new_n517_ = new_n1026_ & new_n1014_ & new_n978_ & new_n966_ & new_n972_ & new_n984_ & new_n1032_ & new_n1020_;
  assign new_n518_ = new_n1026_ & new_n1002_ & new_n978_ & new_n1043_ & new_n1044_ & new_n984_ & new_n1032_ & new_n1008_;
  assign new_n519_ = ~new_n506_;
  assign new_n520_ = ~new_n507_;
  assign new_n521_ = ~new_n508_;
  assign new_n522_ = ~new_n509_;
  assign new_n523_ = ~new_n510_;
  assign new_n524_ = ~new_n511_;
  assign new_n525_ = ~new_n512_;
  assign new_n526_ = ~new_n513_;
  assign new_n527_ = ~new_n516_;
  assign new_n528_ = ~new_n517_;
  assign new_n529_ = ~new_n518_;
  assign new_n530_ = new_n791_ & pi006;
  assign po003 = pi007 & pi006;
  assign new_n532_ = ~new_n530_;
  assign po004 = new_n1489_ | po120 | po094 | po061 | po124 | po054 | po118 | po056 | po095 | po062 | po099;
  assign new_n534_ = pi008 | new_n830_;
  assign po005 = pi009 & new_n534_;
  assign new_n536_ = new_n834_ | new_n899_;
  assign new_n537_ = po065 & new_n536_;
  assign new_n538_ = new_n854_ | new_n537_;
  assign new_n539_ = ~new_n538_;
  assign new_n540_ = new_n874_ | new_n873_;
  assign new_n541_ = new_n520_ | new_n519_;
  assign new_n542_ = new_n522_ | new_n521_;
  assign new_n543_ = new_n524_ | new_n523_;
  assign new_n544_ = new_n526_ | new_n525_;
  assign new_n545_ = new_n541_ & new_n1847_;
  assign new_n546_ = new_n542_ & new_n1848_;
  assign new_n547_ = new_n543_ & new_n1849_;
  assign new_n548_ = pi011 & new_n544_ & pi010;
  assign new_n549_ = new_n545_ | new_n547_ | new_n548_ | new_n546_;
  assign new_n550_ = po160 & po082 & po084 & po083 & new_n552_ & new_n549_;
  assign po006 = new_n1635_ | new_n1636_ | new_n550_;
  assign new_n552_ = ~pi012;
  assign new_n553_ = po160 & pi012;
  assign new_n554_ = po009 | new_n553_;
  assign new_n555_ = new_n1642_ & new_n1640_ & new_n1638_ & new_n1637_ & new_n1639_ & new_n1641_ & new_n588_ & new_n554_ & new_n589_ & new_n584_;
  assign po007 = ~new_n555_;
  assign new_n557_ = ~pi013;
  assign new_n558_ = new_n866_ & new_n863_;
  assign new_n559_ = new_n820_ & new_n862_;
  assign new_n560_ = pi014 & new_n559_;
  assign new_n561_ = ~po165;
  assign new_n562_ = new_n861_ | new_n558_;
  assign new_n563_ = new_n867_ | new_n864_ | new_n657_;
  assign new_n564_ = pi004 & new_n562_;
  assign new_n565_ = pi015 & new_n563_;
  assign new_n566_ = new_n565_ | new_n560_ | new_n564_;
  assign new_n567_ = new_n561_ & new_n566_ & new_n496_;
  assign po008 = ~new_n567_;
  assign new_n569_ = new_n862_ & new_n820_;
  assign new_n570_ = new_n862_ | new_n854_ | new_n843_ | new_n864_ | new_n1715_;
  assign new_n571_ = new_n645_ | pi016 | new_n562_ | new_n569_;
  assign new_n572_ = new_n563_ | new_n1715_;
  assign new_n573_ = po065 & new_n570_;
  assign new_n574_ = pi004 & new_n571_;
  assign new_n575_ = pi015 & new_n572_;
  assign new_n576_ = ~pi017;
  assign new_n577_ = new_n576_ & po052 & new_n496_ & pi018;
  assign new_n578_ = pi019 & new_n1715_;
  assign new_n579_ = new_n1510_ & new_n2007_;
  assign new_n580_ = po065 & new_n579_;
  assign po009 = new_n577_ | new_n574_ | new_n580_ | po160 | new_n560_ | new_n578_ | new_n573_ | new_n575_;
  assign new_n582_ = new_n820_ | po052;
  assign new_n583_ = po065 & new_n582_;
  assign new_n584_ = ~new_n583_;
  assign new_n585_ = ~new_n1677_;
  assign new_n586_ = ~new_n1680_;
  assign new_n587_ = ~new_n1555_;
  assign new_n588_ = ~pi020;
  assign new_n589_ = ~pi021;
  assign po010 = new_n1642_ & new_n1640_ & new_n1638_ & new_n1637_ & new_n1639_ & new_n1641_ & po009 & new_n586_ & new_n495_ & new_n584_ & new_n561_ & new_n585_ & new_n587_ & new_n1719_ & new_n589_ & new_n588_;
  assign new_n591_ = new_n936_ & new_n882_;
  assign new_n592_ = ~new_n591_;
  assign po011 = po047 | po010;
  assign new_n594_ = ~pi022;
  assign new_n595_ = new_n1859_ & new_n2598_;
  assign new_n596_ = new_n1861_ & new_n595_;
  assign new_n597_ = new_n2613_ & new_n595_;
  assign new_n598_ = new_n2613_ & new_n1861_;
  assign new_n599_ = new_n597_ | new_n598_ | new_n596_;
  assign new_n600_ = new_n1847_ & new_n599_;
  assign new_n601_ = new_n2618_ & new_n599_;
  assign new_n602_ = new_n2618_ & new_n1847_;
  assign new_n603_ = new_n601_ | new_n602_ | new_n600_;
  assign new_n604_ = new_n488_ & new_n491_;
  assign new_n605_ = new_n485_ & new_n604_;
  assign new_n606_ = ~new_n491_;
  assign new_n607_ = ~new_n2263_;
  assign new_n608_ = ~new_n2268_;
  assign new_n609_ = new_n607_ & new_n606_;
  assign new_n610_ = new_n608_ & new_n609_;
  assign new_n611_ = new_n2069_ & new_n2258_ & new_n1861_;
  assign new_n612_ = new_n1871_ & new_n2288_ & new_n2070_;
  assign new_n613_ = new_n611_ | new_n612_;
  assign new_n614_ = new_n2071_ & new_n2253_ & new_n1861_;
  assign new_n615_ = new_n1871_ & new_n2283_ & new_n2072_;
  assign new_n616_ = new_n614_ | new_n615_;
  assign new_n617_ = new_n2073_ & new_n2248_ & new_n1861_;
  assign new_n618_ = new_n1871_ & new_n2278_ & new_n2074_;
  assign new_n619_ = new_n617_ | new_n618_;
  assign new_n620_ = new_n2075_ & new_n2233_ & new_n1861_;
  assign new_n621_ = new_n1871_ & new_n606_ & new_n2076_;
  assign new_n622_ = new_n620_ | new_n621_;
  assign new_n623_ = ~new_n622_;
  assign new_n624_ = ~new_n619_;
  assign new_n625_ = ~new_n616_;
  assign new_n626_ = new_n624_ & new_n623_;
  assign new_n627_ = new_n625_ & new_n626_;
  assign new_n628_ = new_n2077_ & new_n2258_ & new_n1859_;
  assign new_n629_ = new_n1870_ & new_n2303_ & new_n2078_;
  assign new_n630_ = new_n628_ | new_n629_;
  assign new_n631_ = new_n2079_ & new_n2253_ & new_n1859_;
  assign new_n632_ = new_n1870_ & new_n2298_ & new_n2080_;
  assign new_n633_ = new_n631_ | new_n632_;
  assign new_n634_ = new_n2081_ & new_n2248_ & new_n1859_;
  assign new_n635_ = new_n1870_ & new_n2293_ & new_n2082_;
  assign new_n636_ = new_n634_ | new_n635_;
  assign new_n637_ = new_n2083_ & new_n2233_ & new_n1859_;
  assign new_n638_ = new_n1870_ & new_n623_ & new_n2084_;
  assign new_n639_ = new_n637_ | new_n638_;
  assign new_n640_ = ~pi023;
  assign new_n641_ = ~new_n1664_;
  assign new_n642_ = new_n641_ & new_n640_;
  assign po012 = ~new_n642_;
  assign new_n644_ = new_n866_ & new_n843_;
  assign new_n645_ = new_n820_ & new_n843_;
  assign new_n646_ = new_n854_ | new_n860_ | new_n644_ | new_n751_ | new_n902_;
  assign new_n647_ = new_n874_ | new_n873_;
  assign new_n648_ = pi004 & new_n646_;
  assign new_n649_ = pi004 & new_n647_;
  assign new_n650_ = new_n645_ & pi015;
  assign po013 = new_n753_ | new_n649_ | new_n650_ | new_n648_;
  assign new_n652_ = ~new_n2308_;
  assign po014 = new_n671_ | pi024;
  assign po015 = new_n672_ & new_n652_;
  assign new_n655_ = pi004 & new_n558_;
  assign new_n656_ = new_n861_ & pi004;
  assign new_n657_ = new_n820_ & new_n863_;
  assign new_n658_ = pi015 & new_n657_;
  assign new_n659_ = new_n862_ & new_n866_ & pi015;
  assign new_n660_ = new_n864_ & pi015;
  assign new_n661_ = ~new_n655_;
  assign new_n662_ = ~new_n656_;
  assign new_n663_ = ~new_n658_;
  assign new_n664_ = ~new_n659_;
  assign new_n665_ = ~new_n660_;
  assign new_n666_ = ~new_n560_;
  assign new_n667_ = new_n665_ & new_n663_ & new_n661_ & new_n662_ & new_n666_ & new_n664_;
  assign new_n668_ = ~new_n667_;
  assign po016 = new_n588_ & new_n496_ & new_n668_ & new_n586_ & new_n589_;
  assign new_n670_ = ~pi020;
  assign new_n671_ = pi025 & new_n670_;
  assign new_n672_ = ~new_n2313_;
  assign new_n673_ = ~new_n2318_;
  assign new_n674_ = pi026 & pi004 & new_n834_;
  assign new_n675_ = new_n1680_ & new_n834_;
  assign new_n676_ = new_n675_ | new_n674_;
  assign po017 = po081 & new_n902_;
  assign po018 = po080 & new_n902_;
  assign po019 = po079 & new_n902_;
  assign po020 = po078 & new_n902_;
  assign po021 = po077 & new_n902_;
  assign po022 = po076 & new_n902_;
  assign po023 = po075 & new_n902_;
  assign po024 = po074 & new_n902_;
  assign po025 = po073 & new_n902_;
  assign po026 = po072 & new_n902_;
  assign po027 = po071 & new_n902_;
  assign po028 = po070 & new_n902_;
  assign new_n689_ = new_n2085_ & new_n2086_ & new_n860_ & pi026 & po065;
  assign new_n690_ = new_n2085_ & new_n2086_ & new_n860_ & pi027 & po065;
  assign new_n691_ = new_n2085_ & new_n2086_ & new_n860_ & pi028 & po065;
  assign new_n692_ = new_n2085_ & new_n2086_ & new_n860_ & pi029 & po065;
  assign new_n693_ = new_n2087_ & new_n2015_ & new_n1884_ & new_n2088_;
  assign po029 = new_n713_ | new_n693_;
  assign new_n695_ = new_n2087_ & new_n2015_ & new_n2888_ & new_n2088_;
  assign po030 = new_n714_ | new_n695_;
  assign new_n697_ = new_n2087_ & new_n2015_ & new_n2883_ & new_n2088_;
  assign po031 = new_n715_ | new_n697_;
  assign new_n699_ = new_n2087_ & new_n2015_ & new_n2878_ & new_n2088_;
  assign po032 = new_n716_ | new_n699_;
  assign new_n701_ = new_n2087_ & new_n2015_ & new_n2873_ & new_n2088_;
  assign po033 = new_n717_ | new_n701_;
  assign new_n703_ = new_n2087_ & new_n2015_ & new_n2868_ & new_n2088_;
  assign po034 = new_n718_ | new_n703_;
  assign new_n705_ = new_n2087_ & new_n2015_ & new_n2863_ & new_n2088_;
  assign po035 = new_n719_ | new_n689_ | new_n705_;
  assign new_n707_ = new_n2087_ & new_n2015_ & new_n2858_ & new_n2088_;
  assign po036 = new_n720_ | new_n690_ | new_n707_;
  assign new_n709_ = new_n2087_ & new_n2015_ & new_n2853_ & new_n2088_;
  assign po037 = new_n721_ | new_n691_ | new_n709_;
  assign new_n711_ = new_n2087_ & new_n2015_ & new_n2848_ & new_n2088_;
  assign po038 = new_n722_ | new_n692_ | new_n711_;
  assign new_n713_ = new_n2090_ & new_n2089_ & new_n902_ & po082 & po065;
  assign new_n714_ = new_n2090_ & new_n2089_ & new_n902_ & po083 & po065;
  assign new_n715_ = new_n2090_ & new_n2089_ & new_n902_ & po084 & po065;
  assign new_n716_ = new_n2090_ & new_n2089_ & new_n902_ & po085 & po065;
  assign new_n717_ = new_n2090_ & new_n2089_ & new_n902_ & po086 & po065;
  assign new_n718_ = new_n2090_ & new_n2089_ & new_n902_ & po087 & po065;
  assign new_n719_ = new_n2090_ & new_n2089_ & new_n902_ & po088 & po065;
  assign new_n720_ = new_n2090_ & new_n2089_ & new_n902_ & po089 & po065;
  assign new_n721_ = new_n2090_ & new_n2089_ & new_n902_ & po090 & po065;
  assign new_n722_ = new_n2090_ & new_n2089_ & new_n902_ & po091 & po065;
  assign new_n723_ = ~pi030;
  assign new_n724_ = ~pi031;
  assign po039 = ~pi032;
  assign new_n726_ = ~new_n499_;
  assign po040 = new_n728_ & new_n726_;
  assign new_n728_ = ~pi033;
  assign new_n729_ = new_n726_ & new_n732_ & pi033;
  assign new_n730_ = new_n726_ & pi034 & new_n728_;
  assign po041 = new_n730_ | new_n729_;
  assign new_n732_ = ~pi034;
  assign new_n733_ = pi033 & pi034;
  assign new_n734_ = new_n726_ & new_n738_ & new_n733_;
  assign new_n735_ = ~new_n733_;
  assign new_n736_ = new_n726_ & pi035 & new_n735_;
  assign po042 = new_n736_ | new_n734_;
  assign new_n738_ = ~pi035;
  assign new_n739_ = new_n733_ & pi035;
  assign new_n740_ = new_n726_ & new_n744_ & new_n739_;
  assign new_n741_ = ~new_n739_;
  assign new_n742_ = new_n726_ & pi036 & new_n741_;
  assign po043 = new_n742_ | new_n740_;
  assign new_n744_ = ~pi036;
  assign new_n745_ = new_n739_ & pi036;
  assign new_n746_ = new_n726_ & new_n750_ & new_n745_;
  assign new_n747_ = ~new_n745_;
  assign new_n748_ = new_n726_ & pi037 & new_n747_;
  assign po044 = new_n748_ | new_n746_;
  assign new_n750_ = ~pi037;
  assign new_n751_ = new_n495_ & new_n872_;
  assign new_n752_ = new_n645_ | new_n751_;
  assign new_n753_ = new_n874_ & pi014;
  assign new_n754_ = po133 & new_n648_ & new_n586_ & new_n496_;
  assign new_n755_ = new_n496_ & new_n752_ & po133 & pi015;
  assign new_n756_ = new_n496_ & new_n874_ & po133 & pi014;
  assign new_n757_ = ~new_n754_;
  assign new_n758_ = ~new_n755_;
  assign new_n759_ = ~new_n756_;
  assign po045 = new_n758_ & new_n759_ & new_n757_;
  assign po046 = new_n673_ & pi038;
  assign new_n762_ = ~new_n673_;
  assign new_n763_ = new_n878_ & pi014;
  assign new_n764_ = ~pi039;
  assign new_n765_ = ~new_n763_;
  assign new_n766_ = po065 & new_n1509_ & new_n1681_;
  assign new_n767_ = new_n1771_ & pi015 & new_n1509_;
  assign new_n768_ = new_n878_ & pi004;
  assign new_n769_ = new_n766_ | pi040 | new_n768_ | new_n767_;
  assign po047 = new_n765_ & new_n769_ & new_n764_;
  assign new_n771_ = pi041 & pi023 & new_n779_;
  assign new_n772_ = pi042 & new_n781_ & new_n779_;
  assign new_n773_ = new_n772_ | new_n771_;
  assign po048 = ~new_n773_;
  assign new_n775_ = ~pi043;
  assign new_n776_ = ~new_n782_;
  assign new_n777_ = new_n640_ & new_n776_ & new_n775_;
  assign new_n778_ = new_n779_ & new_n781_;
  assign new_n779_ = ~new_n777_;
  assign po049 = ~new_n778_;
  assign new_n781_ = ~pi023;
  assign new_n782_ = ~pi042;
  assign new_n783_ = ~pi044;
  assign new_n784_ = pi051 & pi050 & pi049 & pi048 & pi047 & pi045 & pi046;
  assign new_n785_ = pi051 & pi050 & pi049 & pi047 & pi045 & pi046;
  assign new_n786_ = pi051 & pi050 & pi047 & pi045 & pi046;
  assign new_n787_ = pi051 & pi050 & pi045 & pi046;
  assign new_n788_ = pi051 & pi045 & pi046;
  assign new_n789_ = pi045 & pi051;
  assign po050 = ~pi045;
  assign new_n791_ = ~pi007;
  assign new_n792_ = ~pi052;
  assign new_n793_ = ~pi053;
  assign new_n794_ = ~pi054;
  assign new_n795_ = ~pi055;
  assign new_n796_ = ~pi056;
  assign new_n797_ = ~pi029;
  assign new_n798_ = ~pi028;
  assign new_n799_ = ~pi027;
  assign new_n800_ = ~pi026;
  assign new_n801_ = ~pi056;
  assign new_n802_ = ~pi029;
  assign new_n803_ = ~pi028;
  assign new_n804_ = ~pi027;
  assign new_n805_ = ~pi026;
  assign new_n806_ = ~new_n797_;
  assign new_n807_ = ~new_n798_;
  assign new_n808_ = ~new_n799_;
  assign new_n809_ = ~new_n800_;
  assign new_n810_ = ~pi056;
  assign new_n811_ = ~pi029;
  assign new_n812_ = ~pi028;
  assign new_n813_ = ~pi027;
  assign new_n814_ = ~pi026;
  assign new_n815_ = ~new_n796_;
  assign new_n816_ = ~new_n797_;
  assign new_n817_ = ~new_n798_;
  assign new_n818_ = ~new_n799_;
  assign new_n819_ = ~new_n800_;
  assign new_n820_ = new_n1459_ & pi057;
  assign new_n821_ = ~new_n820_;
  assign new_n822_ = ~pi058;
  assign new_n823_ = ~pi059;
  assign new_n824_ = ~pi060;
  assign new_n825_ = ~pi061;
  assign new_n826_ = ~pi062;
  assign new_n827_ = ~pi063;
  assign new_n828_ = pi064 & new_n823_ & pi058;
  assign new_n829_ = pi063 & new_n1781_ & new_n828_;
  assign new_n830_ = pi059 & new_n822_ & pi009 & pi064;
  assign new_n831_ = new_n827_ & new_n828_;
  assign new_n832_ = ~new_n831_;
  assign new_n833_ = new_n794_ & new_n795_ & new_n793_;
  assign new_n834_ = new_n793_ & new_n794_ & pi055;
  assign new_n835_ = new_n793_ & new_n795_ & pi054;
  assign new_n836_ = pi055 & new_n794_ & pi053;
  assign new_n837_ = pi054 & pi055 & pi053;
  assign new_n838_ = ~pi055;
  assign new_n839_ = pi054 & new_n838_ & pi053;
  assign po051 = new_n796_ & new_n899_;
  assign new_n841_ = ~pi065;
  assign new_n842_ = ~pi066;
  assign new_n843_ = pi056 & new_n899_;
  assign new_n844_ = pi029 & new_n798_ & po051;
  assign new_n845_ = pi029 & pi028 & po051;
  assign new_n846_ = pi066 & new_n841_ & po051 & new_n798_ & new_n797_;
  assign new_n847_ = new_n842_ & pi065 & po051 & new_n798_ & new_n797_;
  assign new_n848_ = pi066 & pi065 & po051 & new_n798_ & new_n797_;
  assign new_n849_ = new_n842_ & new_n841_ & pi028 & new_n899_ & new_n797_ & new_n796_;
  assign new_n850_ = pi066 & new_n841_ & pi028 & new_n899_ & new_n797_ & new_n796_;
  assign new_n851_ = new_n842_ & pi065 & pi028 & new_n899_ & new_n797_ & new_n796_;
  assign new_n852_ = new_n842_ & new_n841_ & po051 & new_n798_ & new_n797_;
  assign new_n853_ = pi066 & pi065 & pi028 & new_n899_ & new_n797_ & new_n796_;
  assign new_n854_ = pi056 & new_n834_;
  assign new_n855_ = new_n797_ & new_n834_ & new_n798_ & new_n796_;
  assign new_n856_ = new_n797_ & new_n834_ & pi028 & new_n796_;
  assign new_n857_ = pi029 & new_n834_ & new_n798_ & new_n796_;
  assign new_n858_ = new_n796_ & pi055 & pi054 & pi029 & new_n793_;
  assign new_n859_ = new_n796_ & pi055 & pi054 & new_n797_ & new_n793_;
  assign new_n860_ = new_n793_ & pi054 & pi056 & pi055;
  assign new_n861_ = pi029 & new_n834_ & pi028 & new_n796_;
  assign new_n862_ = new_n847_ | new_n845_ | new_n851_ | new_n849_ | new_n848_ | new_n850_ | new_n844_ | new_n846_;
  assign new_n863_ = new_n853_ | new_n852_;
  assign new_n864_ = new_n856_ | new_n857_ | new_n855_;
  assign new_n865_ = ~new_n820_;
  assign new_n866_ = new_n821_ | new_n865_;
  assign new_n867_ = new_n862_ & new_n866_;
  assign new_n868_ = new_n804_ & new_n802_ & new_n835_ & new_n801_ & new_n809_ & new_n803_;
  assign new_n869_ = new_n808_ & new_n802_ & new_n835_ & new_n801_ & new_n805_ & new_n803_;
  assign new_n870_ = new_n808_ & new_n802_ & new_n835_ & new_n801_ & new_n809_ & new_n803_;
  assign new_n871_ = new_n804_ & new_n802_ & new_n835_ & new_n801_ & new_n805_ & new_n807_;
  assign new_n872_ = new_n804_ & new_n802_ & new_n835_ & new_n801_ & new_n809_ & new_n807_;
  assign new_n873_ = new_n808_ & new_n802_ & new_n835_ & new_n801_ & new_n805_ & new_n807_;
  assign new_n874_ = new_n808_ & new_n802_ & new_n835_ & new_n801_ & new_n809_ & new_n807_;
  assign new_n875_ = new_n804_ & new_n806_ & new_n835_ & new_n801_ & new_n805_ & new_n803_;
  assign new_n876_ = new_n813_ & new_n816_ & new_n835_ & new_n810_ & new_n819_ & new_n812_;
  assign new_n877_ = new_n818_ & new_n816_ & new_n835_ & new_n810_ & new_n814_ & new_n812_;
  assign new_n878_ = new_n818_ & new_n816_ & new_n835_ & new_n810_ & new_n819_ & new_n812_;
  assign new_n879_ = new_n813_ & new_n816_ & new_n835_ & new_n810_ & new_n819_ & new_n817_;
  assign new_n880_ = new_n818_ & new_n816_ & new_n835_ & new_n810_ & new_n814_ & new_n817_;
  assign new_n881_ = new_n818_ & new_n816_ & new_n835_ & new_n810_ & new_n819_ & new_n817_;
  assign new_n882_ = new_n813_ & new_n811_ & new_n835_ & new_n815_ & new_n814_ & new_n812_;
  assign new_n883_ = new_n813_ & new_n811_ & new_n835_ & new_n815_ & new_n819_ & new_n812_;
  assign new_n884_ = new_n818_ & new_n811_ & new_n835_ & new_n815_ & new_n814_ & new_n812_;
  assign new_n885_ = ~new_n883_;
  assign new_n886_ = ~new_n884_;
  assign new_n887_ = ~new_n882_;
  assign new_n888_ = new_n886_ & new_n815_ & new_n835_ & new_n887_ & new_n885_;
  assign new_n889_ = new_n813_ & new_n811_ & new_n835_ & new_n810_ & new_n814_ & new_n812_;
  assign new_n890_ = new_n813_ & new_n817_ & new_n835_ & new_n816_ & new_n814_ & new_n810_;
  assign new_n891_ = new_n889_ | new_n890_ | new_n888_;
  assign new_n892_ = new_n881_ | new_n880_;
  assign new_n893_ = ~pi067;
  assign new_n894_ = new_n501_ & new_n893_ & new_n892_;
  assign new_n895_ = new_n894_ | new_n858_ | new_n833_;
  assign po052 = new_n1653_ & new_n1651_ & new_n1652_ & pi068 & new_n895_;
  assign new_n897_ = ~po052;
  assign new_n898_ = ~pi016;
  assign new_n899_ = new_n833_ & new_n898_;
  assign new_n900_ = new_n880_ & new_n898_;
  assign new_n901_ = new_n881_ & new_n898_;
  assign new_n902_ = new_n858_ & new_n898_;
  assign new_n903_ = ~new_n891_;
  assign new_n904_ = ~new_n836_;
  assign new_n905_ = ~new_n839_;
  assign new_n906_ = ~new_n837_;
  assign new_n907_ = new_n905_ & new_n903_ & new_n906_ & new_n904_;
  assign po053 = new_n641_ & new_n1049_ & po052 & pi019 & new_n1708_;
  assign new_n909_ = new_n898_ & new_n503_;
  assign new_n910_ = new_n909_ | pi069;
  assign po054 = pi070 & pi052;
  assign po055 = new_n530_ & pi071;
  assign po056 = pi052 & pi071;
  assign po057 = pi071 & new_n910_ & pi072;
  assign po058 = new_n530_ & pi031;
  assign po059 = pi070 & pi073;
  assign po060 = pi031 & pi073;
  assign new_n918_ = ~new_n724_;
  assign new_n919_ = ~new_n792_;
  assign po061 = new_n919_ & new_n918_;
  assign new_n921_ = pi007 | new_n1629_;
  assign po062 = pi074 & pi052 & new_n921_;
  assign new_n923_ = po186 & new_n891_;
  assign new_n924_ = ~new_n923_;
  assign new_n925_ = ~new_n907_;
  assign new_n926_ = ~new_n1715_;
  assign new_n927_ = new_n925_ & new_n926_ & new_n924_;
  assign new_n928_ = ~new_n927_;
  assign new_n929_ = ~new_n950_;
  assign new_n930_ = new_n929_ & new_n641_ & new_n928_;
  assign po063 = ~new_n930_;
  assign new_n932_ = new_n826_ & new_n824_ & pi075 & pi019 & new_n825_;
  assign new_n933_ = ~new_n892_;
  assign po064 = new_n933_ & new_n932_;
  assign po065 = pi069 | pi076;
  assign new_n936_ = ~po065;
  assign new_n937_ = ~new_n873_;
  assign new_n938_ = ~new_n872_;
  assign new_n939_ = new_n938_ & new_n937_;
  assign new_n940_ = new_n831_ | new_n1998_ | new_n829_ | pi039;
  assign new_n941_ = pi077 & new_n874_;
  assign new_n942_ = ~new_n939_;
  assign new_n943_ = ~new_n1359_;
  assign new_n944_ = new_n943_ & new_n942_;
  assign new_n945_ = new_n944_ | new_n1066_ | new_n941_;
  assign new_n946_ = new_n830_ | new_n940_;
  assign new_n947_ = new_n1780_ & new_n832_ & new_n945_;
  assign new_n948_ = new_n1771_ & new_n946_;
  assign new_n949_ = new_n496_ & pi078;
  assign new_n950_ = pi005 | new_n947_ | new_n949_ | pi039 | new_n829_ | new_n948_ | pi021;
  assign new_n951_ = pi028 & new_n498_;
  assign new_n952_ = ~new_n498_;
  assign new_n953_ = new_n955_ & new_n952_;
  assign po066 = new_n953_ | new_n951_;
  assign new_n955_ = ~pi079;
  assign new_n956_ = pi029 & new_n498_;
  assign new_n957_ = new_n960_ & new_n953_;
  assign new_n958_ = pi079 & pi080 & new_n952_;
  assign po067 = new_n957_ | new_n958_ | new_n956_;
  assign new_n960_ = ~pi080;
  assign new_n961_ = ~new_n2358_;
  assign new_n962_ = ~new_n2363_;
  assign new_n963_ = ~new_n2368_;
  assign new_n964_ = ~new_n2373_;
  assign new_n965_ = new_n1864_ & new_n963_ & new_n961_ & new_n962_ & new_n592_ & new_n964_;
  assign new_n966_ = ~new_n965_;
  assign new_n967_ = ~new_n2378_;
  assign new_n968_ = ~new_n2383_;
  assign new_n969_ = ~new_n2388_;
  assign new_n970_ = ~new_n2393_;
  assign new_n971_ = pi081 & new_n969_ & new_n967_ & new_n968_ & new_n592_ & new_n970_;
  assign new_n972_ = ~new_n971_;
  assign new_n973_ = ~new_n2398_;
  assign new_n974_ = ~new_n2403_;
  assign new_n975_ = ~new_n2408_;
  assign new_n976_ = ~new_n2413_;
  assign new_n977_ = new_n1849_ & new_n975_ & new_n973_ & new_n974_ & new_n592_ & new_n976_;
  assign new_n978_ = ~new_n977_;
  assign new_n979_ = ~new_n2418_;
  assign new_n980_ = ~new_n2423_;
  assign new_n981_ = ~new_n2428_;
  assign new_n982_ = ~new_n2433_;
  assign new_n983_ = new_n1849_ & new_n981_ & new_n979_ & new_n980_ & new_n592_ & new_n982_;
  assign new_n984_ = ~new_n983_;
  assign new_n985_ = ~new_n2438_;
  assign new_n986_ = ~new_n2443_;
  assign new_n987_ = ~new_n2448_;
  assign new_n988_ = ~new_n2453_;
  assign new_n989_ = new_n1863_ & new_n987_ & new_n985_ & new_n986_ & new_n592_ & new_n988_;
  assign new_n990_ = ~new_n989_;
  assign new_n991_ = ~new_n2458_;
  assign new_n992_ = ~new_n2463_;
  assign new_n993_ = ~new_n2468_;
  assign new_n994_ = ~new_n2473_;
  assign new_n995_ = pi082 & new_n993_ & new_n991_ & new_n992_ & new_n592_ & new_n994_;
  assign new_n996_ = ~new_n995_;
  assign new_n997_ = ~new_n2478_;
  assign new_n998_ = ~new_n2483_;
  assign new_n999_ = ~new_n2488_;
  assign new_n1000_ = ~new_n2493_;
  assign new_n1001_ = new_n1848_ & new_n999_ & new_n997_ & new_n998_ & new_n592_ & new_n1000_;
  assign new_n1002_ = ~new_n1001_;
  assign new_n1003_ = ~new_n2498_;
  assign new_n1004_ = ~new_n2503_;
  assign new_n1005_ = ~new_n2508_;
  assign new_n1006_ = ~new_n2513_;
  assign new_n1007_ = new_n1848_ & new_n1005_ & new_n1003_ & new_n1004_ & new_n592_ & new_n1006_;
  assign new_n1008_ = ~new_n1007_;
  assign new_n1009_ = ~new_n2518_;
  assign new_n1010_ = ~new_n2523_;
  assign new_n1011_ = ~new_n2528_;
  assign new_n1012_ = ~new_n2533_;
  assign new_n1013_ = new_n1862_ & new_n1011_ & new_n1009_ & new_n1010_ & new_n592_ & new_n1012_;
  assign new_n1014_ = ~new_n1013_;
  assign new_n1015_ = ~new_n2538_;
  assign new_n1016_ = ~new_n2543_;
  assign new_n1017_ = ~new_n2548_;
  assign new_n1018_ = ~new_n2553_;
  assign new_n1019_ = pi083 & new_n1017_ & new_n1015_ & new_n1016_ & new_n592_ & new_n1018_;
  assign new_n1020_ = ~new_n1019_;
  assign new_n1021_ = ~new_n2558_;
  assign new_n1022_ = ~new_n2563_;
  assign new_n1023_ = ~new_n2568_;
  assign new_n1024_ = ~new_n2573_;
  assign new_n1025_ = new_n1847_ & new_n1023_ & new_n1021_ & new_n1022_ & new_n592_ & new_n1024_;
  assign new_n1026_ = ~new_n1025_;
  assign new_n1027_ = ~new_n2578_;
  assign new_n1028_ = ~new_n2583_;
  assign new_n1029_ = ~new_n2588_;
  assign new_n1030_ = ~new_n2593_;
  assign new_n1031_ = new_n1847_ & new_n1029_ & new_n1027_ & new_n1028_ & new_n592_ & new_n1030_;
  assign new_n1032_ = ~new_n1031_;
  assign new_n1033_ = ~new_n1339_;
  assign new_n1034_ = ~new_n1337_;
  assign new_n1035_ = ~new_n1335_;
  assign new_n1036_ = ~new_n1333_;
  assign new_n1037_ = new_n1865_ & new_n1035_ & new_n1033_ & new_n1034_ & new_n592_ & new_n1036_;
  assign new_n1038_ = pi010 & new_n1035_ & new_n1033_ & new_n1034_ & new_n592_ & new_n1333_;
  assign new_n1039_ = pi011 & pi010 & new_n1036_ & new_n1033_ & new_n1034_ & new_n592_ & new_n1335_;
  assign new_n1040_ = pi011 & pi010 & new_n1333_ & new_n1335_ & new_n1033_ & new_n592_ & new_n1034_;
  assign new_n1041_ = ~new_n1037_;
  assign new_n1042_ = ~new_n1038_;
  assign new_n1043_ = ~new_n1039_;
  assign new_n1044_ = ~new_n1040_;
  assign new_n1045_ = po065 & new_n928_;
  assign new_n1046_ = new_n910_ & new_n892_ & pi004 & po052;
  assign new_n1047_ = pi004 & new_n891_;
  assign new_n1048_ = new_n932_ & new_n892_;
  assign new_n1049_ = ~new_n940_;
  assign new_n1050_ = new_n1045_ | new_n1047_ | new_n1048_ | new_n1046_;
  assign po068 = new_n641_ & new_n1050_ & new_n1049_;
  assign new_n1052_ = ~pi004;
  assign new_n1053_ = pi084 & new_n1532_ & new_n1524_ & new_n1072_ & new_n1715_;
  assign new_n1054_ = ~new_n1053_;
  assign new_n1055_ = ~new_n869_;
  assign new_n1056_ = ~new_n875_;
  assign new_n1057_ = ~new_n876_;
  assign new_n1058_ = ~new_n877_;
  assign new_n1059_ = ~new_n868_;
  assign new_n1060_ = ~new_n879_;
  assign new_n1061_ = new_n1059_ & new_n1057_ & new_n1055_ & new_n1054_ & new_n1056_ & new_n1060_ & new_n1058_;
  assign new_n1062_ = ~new_n1046_;
  assign new_n1063_ = new_n1062_ & new_n1061_ & pi004 & new_n903_;
  assign new_n1064_ = ~new_n1061_;
  assign new_n1065_ = ~new_n1052_;
  assign new_n1066_ = new_n1065_ & new_n1064_;
  assign new_n1067_ = new_n644_ | new_n854_ | new_n2007_;
  assign new_n1068_ = pi015 & new_n1067_;
  assign new_n1069_ = pi014 & new_n1715_;
  assign new_n1070_ = new_n1068_ | new_n1069_ | new_n1063_;
  assign po069 = new_n641_ & new_n1070_ & new_n1049_;
  assign new_n1072_ = ~pi015;
  assign new_n1073_ = new_n2091_ & pi085 & new_n1459_;
  assign new_n1074_ = new_n2091_ & pi086 & new_n1459_;
  assign new_n1075_ = new_n2091_ & pi087 & new_n1459_;
  assign new_n1076_ = new_n2091_ & pi088 & new_n1459_;
  assign new_n1077_ = new_n2091_ & pi089 & new_n1459_;
  assign new_n1078_ = new_n2091_ & pi090 & new_n1459_;
  assign new_n1079_ = new_n2091_ & pi091 & new_n1459_;
  assign new_n1080_ = new_n2091_ & pi092 & new_n1459_;
  assign new_n1081_ = new_n2091_ & pi093 & new_n1459_;
  assign new_n1082_ = new_n2091_ & pi094 & new_n1459_;
  assign new_n1083_ = new_n2091_ & pi095 & new_n1459_;
  assign new_n1084_ = new_n2091_ & pi096 & new_n1459_;
  assign new_n1085_ = new_n2007_ & pi097 & new_n2092_;
  assign new_n1086_ = new_n1073_ | new_n1085_;
  assign new_n1087_ = new_n2007_ & pi098 & new_n2092_;
  assign new_n1088_ = new_n1074_ | new_n1087_;
  assign new_n1089_ = new_n2007_ & pi099 & new_n2092_;
  assign new_n1090_ = new_n1075_ | new_n1089_;
  assign new_n1091_ = new_n2007_ & pi100 & new_n2092_;
  assign new_n1092_ = new_n1076_ | new_n1091_;
  assign new_n1093_ = new_n2007_ & pi101 & new_n2092_;
  assign new_n1094_ = new_n1077_ | new_n1093_;
  assign new_n1095_ = new_n2007_ & pi102 & new_n2092_;
  assign new_n1096_ = new_n1078_ | new_n1095_;
  assign new_n1097_ = new_n2007_ & pi103 & new_n2092_;
  assign new_n1098_ = new_n1079_ | new_n1097_;
  assign new_n1099_ = new_n2007_ & pi104 & new_n2092_;
  assign new_n1100_ = new_n1080_ | new_n1099_;
  assign new_n1101_ = new_n2007_ & pi105 & new_n2092_;
  assign new_n1102_ = new_n1081_ | new_n1101_;
  assign new_n1103_ = new_n2007_ & pi106 & new_n2092_;
  assign new_n1104_ = new_n1082_ | new_n1103_;
  assign new_n1105_ = new_n2007_ & pi107 & new_n2092_;
  assign new_n1106_ = new_n1083_ | new_n1105_;
  assign new_n1107_ = new_n2007_ & pi108 & new_n2092_;
  assign new_n1108_ = new_n1084_ | new_n1107_;
  assign new_n1109_ = new_n2093_ & pi109 & new_n1459_;
  assign new_n1110_ = new_n2093_ & pi110 & new_n1459_;
  assign new_n1111_ = new_n2093_ & pi111 & new_n1459_;
  assign new_n1112_ = new_n2093_ & pi112 & new_n1459_;
  assign new_n1113_ = new_n2093_ & pi113 & new_n1459_;
  assign new_n1114_ = new_n2093_ & pi114 & new_n1459_;
  assign new_n1115_ = new_n2093_ & pi115 & new_n1459_;
  assign new_n1116_ = new_n2093_ & pi116 & new_n1459_;
  assign new_n1117_ = new_n2093_ & pi117 & new_n1459_;
  assign new_n1118_ = new_n2093_ & pi118 & new_n1459_;
  assign new_n1119_ = new_n2007_ & pi119 & new_n2094_;
  assign new_n1120_ = new_n1109_ | new_n1119_;
  assign new_n1121_ = new_n2007_ & pi120 & new_n2094_;
  assign new_n1122_ = new_n1110_ | new_n1121_;
  assign new_n1123_ = new_n2007_ & pi121 & new_n2094_;
  assign new_n1124_ = new_n1111_ | new_n1123_;
  assign new_n1125_ = new_n2007_ & pi122 & new_n2094_;
  assign new_n1126_ = new_n1112_ | new_n1125_;
  assign new_n1127_ = new_n2007_ & pi123 & new_n2094_;
  assign new_n1128_ = new_n1113_ | new_n1127_;
  assign new_n1129_ = new_n2007_ & pi124 & new_n2094_;
  assign new_n1130_ = new_n1114_ | new_n1129_;
  assign new_n1131_ = new_n2007_ & pi125 & new_n2094_;
  assign new_n1132_ = new_n1115_ | new_n1131_;
  assign new_n1133_ = new_n2007_ & pi126 & new_n2094_;
  assign new_n1134_ = new_n1116_ | new_n1133_;
  assign new_n1135_ = new_n2007_ & pi127 & new_n2094_;
  assign new_n1136_ = new_n1117_ | new_n1135_;
  assign new_n1137_ = new_n2007_ & pi128 & new_n2094_;
  assign new_n1138_ = new_n1118_ | new_n1137_;
  assign new_n1139_ = new_n2095_ & new_n2096_ & pi051 & new_n1715_;
  assign new_n1140_ = new_n2095_ & new_n2096_ & pi046 & new_n1715_;
  assign new_n1141_ = new_n2095_ & new_n2096_ & pi050 & new_n1715_;
  assign new_n1142_ = new_n2095_ & new_n2096_ & pi047 & new_n1715_;
  assign new_n1143_ = new_n2095_ & new_n2096_ & pi049 & new_n1715_;
  assign new_n1144_ = new_n2095_ & new_n2096_ & pi048 & new_n1715_;
  assign new_n1145_ = new_n2095_ & new_n2096_ & pi129 & new_n1715_;
  assign new_n1146_ = new_n2095_ & new_n2096_ & pi051 & new_n1715_;
  assign new_n1147_ = new_n1139_ | new_n1155_;
  assign new_n1148_ = new_n1140_ | new_n1156_;
  assign new_n1149_ = new_n1141_ | new_n1157_;
  assign new_n1150_ = new_n1142_ | new_n1158_;
  assign new_n1151_ = new_n1143_ | new_n1159_;
  assign new_n1152_ = new_n1144_ | new_n1160_;
  assign new_n1153_ = new_n1145_ | new_n1161_;
  assign new_n1154_ = new_n1146_ | new_n1162_;
  assign new_n1155_ = new_n1485_ & new_n2097_ & new_n1086_ & new_n2098_;
  assign new_n1156_ = new_n1485_ & new_n2097_ & new_n1088_ & new_n2098_;
  assign new_n1157_ = new_n1485_ & new_n2097_ & new_n1090_ & new_n2098_;
  assign new_n1158_ = new_n1485_ & new_n2097_ & new_n1092_ & new_n2098_;
  assign new_n1159_ = new_n1485_ & new_n2097_ & new_n1094_ & new_n2098_;
  assign new_n1160_ = new_n1485_ & new_n2097_ & new_n1096_ & new_n2098_;
  assign new_n1161_ = new_n1485_ & new_n2097_ & new_n1098_ & new_n2098_;
  assign new_n1162_ = new_n1485_ & new_n2097_ & new_n1100_ & new_n2098_;
  assign new_n1163_ = new_n2099_ & new_n2100_ & pi045 & new_n1715_;
  assign new_n1164_ = new_n2101_ & new_n2102_ & new_n860_ & new_n1510_ & pi026 & new_n1072_;
  assign new_n1165_ = new_n1172_ | new_n1164_;
  assign new_n1166_ = new_n2101_ & new_n2102_ & new_n860_ & new_n1510_ & pi027 & new_n1072_;
  assign new_n1167_ = new_n1173_ | new_n1166_;
  assign new_n1168_ = new_n2101_ & new_n2102_ & new_n860_ & new_n1510_ & pi028 & new_n1072_;
  assign new_n1169_ = new_n1174_ | new_n1168_;
  assign new_n1170_ = new_n2101_ & new_n2102_ & new_n860_ & new_n1510_ & pi029 & new_n1072_;
  assign new_n1171_ = new_n1175_ | new_n1163_ | new_n1170_;
  assign new_n1172_ = new_n1485_ & new_n2103_ & new_n1132_ & new_n2104_;
  assign new_n1173_ = new_n1485_ & new_n2103_ & new_n1134_ & new_n2104_;
  assign new_n1174_ = new_n1485_ & new_n2103_ & new_n1136_ & new_n2104_;
  assign new_n1175_ = new_n1485_ & new_n2103_ & new_n1138_ & new_n2104_;
  assign new_n1176_ = new_n2106_ & pi130;
  assign new_n1177_ = new_n2106_ & pi131;
  assign new_n1178_ = new_n2106_ & pi132;
  assign new_n1179_ = new_n2106_ & pi133;
  assign new_n1180_ = new_n2106_ & pi134;
  assign new_n1181_ = new_n2106_ & pi003;
  assign new_n1182_ = new_n2106_ & pi002;
  assign new_n1183_ = new_n2106_ & pi001;
  assign new_n1184_ = new_n2106_ & pi000;
  assign new_n1185_ = new_n1472_ & pi135 & new_n2107_;
  assign new_n1186_ = new_n1176_ | new_n1185_;
  assign new_n1187_ = new_n1472_ & pi136 & new_n2107_;
  assign new_n1188_ = new_n1177_ | new_n1187_;
  assign new_n1189_ = new_n1472_ & pi137 & new_n2107_;
  assign new_n1190_ = new_n1178_ | new_n1189_;
  assign new_n1191_ = new_n1472_ & pi130 & new_n2107_;
  assign new_n1192_ = new_n1179_ | new_n1191_;
  assign new_n1193_ = new_n1472_ & pi131 & new_n2107_;
  assign new_n1194_ = new_n1180_ | new_n1193_;
  assign new_n1195_ = new_n1472_ & pi132 & new_n2107_;
  assign new_n1196_ = new_n1181_ | new_n1195_;
  assign new_n1197_ = new_n1472_ & pi133 & new_n2107_;
  assign new_n1198_ = new_n1182_ | new_n1197_;
  assign new_n1199_ = new_n1472_ & pi134 & new_n2107_;
  assign new_n1200_ = new_n1183_ | new_n1199_;
  assign new_n1201_ = new_n1472_ & pi003 & new_n2107_;
  assign new_n1202_ = new_n1184_ | new_n1201_;
  assign new_n1203_ = new_n1472_ & pi002 & new_n2107_;
  assign new_n1204_ = new_n2106_ | new_n1203_;
  assign new_n1205_ = new_n1472_ & pi001 & new_n2107_;
  assign new_n1206_ = new_n2106_ | new_n1205_;
  assign new_n1207_ = new_n1472_ & pi000 & new_n2107_;
  assign new_n1208_ = new_n2106_ | new_n1207_;
  assign new_n1209_ = new_n1719_ & po052;
  assign new_n1210_ = ~new_n1209_;
  assign new_n1211_ = new_n2108_ & new_n1147_ & new_n1210_;
  assign new_n1212_ = new_n2108_ & new_n1148_ & new_n1210_;
  assign new_n1213_ = new_n2108_ & new_n1149_ & new_n1210_;
  assign new_n1214_ = new_n2108_ & new_n1150_ & new_n1210_;
  assign new_n1215_ = new_n2108_ & new_n1151_ & new_n1210_;
  assign new_n1216_ = new_n2108_ & new_n1152_ & new_n1210_;
  assign new_n1217_ = new_n2108_ & new_n1153_ & new_n1210_;
  assign new_n1218_ = new_n1209_ & new_n1200_ & new_n2109_;
  assign new_n1219_ = new_n1211_ | new_n1218_;
  assign new_n1220_ = new_n1209_ & new_n1202_ & new_n2109_;
  assign new_n1221_ = new_n1212_ | new_n1220_;
  assign new_n1222_ = new_n1209_ & new_n1204_ & new_n2109_;
  assign new_n1223_ = new_n1213_ | new_n1222_;
  assign new_n1224_ = new_n1209_ & new_n1206_ & new_n2109_;
  assign new_n1225_ = new_n1214_ | new_n1224_;
  assign new_n1226_ = new_n1209_ & new_n1208_ & new_n2109_;
  assign new_n1227_ = new_n1215_ | new_n1226_;
  assign new_n1228_ = new_n1209_ & new_n2106_ & new_n2109_;
  assign new_n1229_ = new_n1216_ | new_n1228_;
  assign new_n1230_ = new_n1209_ & new_n2109_ & new_n1472_ & new_n2107_;
  assign new_n1231_ = new_n1217_ | new_n1230_;
  assign new_n1232_ = new_n2110_ & new_n1210_ & new_n2103_ & new_n2104_ & new_n1485_ & new_n1120_;
  assign new_n1233_ = new_n2110_ & new_n1210_ & new_n2103_ & new_n2104_ & new_n1485_ & new_n1122_;
  assign new_n1234_ = new_n2110_ & new_n1210_ & new_n2103_ & new_n2104_ & new_n1485_ & new_n1124_;
  assign new_n1235_ = new_n2110_ & new_n1210_ & new_n2103_ & new_n2104_ & new_n1485_ & new_n1126_;
  assign new_n1236_ = new_n2110_ & new_n1210_ & new_n2103_ & new_n2104_ & new_n1485_ & new_n1128_;
  assign new_n1237_ = new_n2110_ & new_n1210_ & new_n2103_ & new_n2104_ & new_n1485_ & new_n1130_;
  assign new_n1238_ = new_n2110_ & new_n1165_ & new_n1210_;
  assign new_n1239_ = new_n2110_ & new_n1167_ & new_n1210_;
  assign new_n1240_ = new_n2110_ & new_n1169_ & new_n1210_;
  assign new_n1241_ = new_n2110_ & new_n1171_ & new_n1210_;
  assign new_n1242_ = new_n1209_ & new_n2111_ & new_n2106_ & pi135;
  assign new_n1243_ = new_n1232_ | new_n1242_;
  assign new_n1244_ = new_n1209_ & new_n2111_ & new_n2106_ & pi136;
  assign new_n1245_ = new_n1233_ | new_n1244_;
  assign new_n1246_ = new_n1209_ & new_n2111_ & new_n2106_ & pi137;
  assign new_n1247_ = new_n1234_ | new_n1246_;
  assign new_n1248_ = new_n1209_ & new_n1186_ & new_n2111_;
  assign new_n1249_ = new_n1235_ | new_n1248_;
  assign new_n1250_ = new_n1209_ & new_n1188_ & new_n2111_;
  assign new_n1251_ = new_n1236_ | new_n1250_;
  assign new_n1252_ = new_n1209_ & new_n1190_ & new_n2111_;
  assign new_n1253_ = new_n1237_ | new_n1252_;
  assign new_n1254_ = new_n1209_ & new_n1192_ & new_n2111_;
  assign new_n1255_ = new_n1238_ | new_n1254_;
  assign new_n1256_ = new_n1209_ & new_n1194_ & new_n2111_;
  assign new_n1257_ = new_n1239_ | new_n1256_;
  assign new_n1258_ = new_n1209_ & new_n1196_ & new_n2111_;
  assign new_n1259_ = new_n1240_ | new_n1258_;
  assign new_n1260_ = new_n1209_ & new_n1198_ & new_n2111_;
  assign new_n1261_ = new_n1241_ | new_n1260_;
  assign new_n1262_ = new_n2112_ & new_n1219_ & new_n1486_;
  assign new_n1263_ = new_n2112_ & new_n1221_ & new_n1486_;
  assign new_n1264_ = new_n2112_ & new_n1223_ & new_n1486_;
  assign new_n1265_ = new_n2112_ & new_n1225_ & new_n1486_;
  assign new_n1266_ = new_n2112_ & new_n1227_ & new_n1486_;
  assign new_n1267_ = new_n2112_ & new_n1229_ & new_n1486_;
  assign new_n1268_ = new_n2112_ & new_n1231_ & new_n1486_;
  assign new_n1269_ = new_n2112_ & new_n1486_ & new_n1210_ & new_n2108_ & new_n1154_;
  assign new_n1270_ = new_n2112_ & new_n1486_ & new_n1210_ & new_n2097_ & new_n2098_ & new_n1102_ & new_n2108_ & new_n1485_;
  assign new_n1271_ = new_n2112_ & new_n1486_ & new_n1210_ & new_n2097_ & new_n2098_ & new_n1104_ & new_n2108_ & new_n1485_;
  assign new_n1272_ = new_n2112_ & new_n1486_ & new_n1210_ & new_n2097_ & new_n2098_ & new_n1106_ & new_n2108_ & new_n1485_;
  assign new_n1273_ = new_n2112_ & new_n1486_ & new_n1210_ & new_n2097_ & new_n2098_ & new_n1108_ & new_n2108_ & new_n1485_;
  assign new_n1274_ = new_n1481_ & pi135 & new_n2113_;
  assign po070 = new_n1262_ | new_n1274_;
  assign new_n1276_ = new_n1481_ & pi136 & new_n2113_;
  assign po071 = new_n1263_ | new_n1276_;
  assign new_n1278_ = new_n1481_ & pi137 & new_n2113_;
  assign po072 = new_n1264_ | new_n1278_;
  assign new_n1280_ = new_n1481_ & pi130 & new_n2113_;
  assign po073 = new_n1265_ | new_n1280_;
  assign new_n1282_ = new_n1481_ & pi131 & new_n2113_;
  assign po074 = new_n1266_ | new_n1282_;
  assign new_n1284_ = new_n1481_ & pi132 & new_n2113_;
  assign po075 = new_n1267_ | new_n1284_;
  assign new_n1286_ = new_n1481_ & pi133 & new_n2113_;
  assign po076 = new_n1268_ | new_n1286_;
  assign new_n1288_ = new_n1481_ & pi134 & new_n2113_;
  assign po077 = new_n1269_ | new_n1288_;
  assign new_n1290_ = new_n1481_ & pi003 & new_n2113_;
  assign po078 = new_n1270_ | new_n1290_;
  assign new_n1292_ = new_n1481_ & pi002 & new_n2113_;
  assign po079 = new_n1271_ | new_n1292_;
  assign new_n1294_ = new_n1481_ & pi001 & new_n2113_;
  assign po080 = new_n1272_ | new_n1294_;
  assign new_n1296_ = new_n1481_ & pi000 & new_n2113_;
  assign po081 = new_n1273_ | new_n1296_;
  assign new_n1298_ = new_n2114_ & new_n1243_ & new_n1486_;
  assign new_n1299_ = new_n2114_ & new_n1245_ & new_n1486_;
  assign new_n1300_ = new_n2114_ & new_n1247_ & new_n1486_;
  assign new_n1301_ = new_n2114_ & new_n1249_ & new_n1486_;
  assign new_n1302_ = new_n2114_ & new_n1251_ & new_n1486_;
  assign new_n1303_ = new_n2114_ & new_n1253_ & new_n1486_;
  assign new_n1304_ = new_n2114_ & new_n1255_ & new_n1486_;
  assign new_n1305_ = new_n2114_ & new_n1257_ & new_n1486_;
  assign new_n1306_ = new_n2114_ & new_n1259_ & new_n1486_;
  assign new_n1307_ = new_n2114_ & new_n1261_ & new_n1486_;
  assign new_n1308_ = new_n1481_ & pi138 & new_n2115_;
  assign po082 = new_n1298_ | new_n1308_;
  assign new_n1310_ = new_n1481_ & pi139 & new_n2115_;
  assign po083 = new_n1299_ | new_n1310_;
  assign new_n1312_ = new_n1481_ & pi140 & new_n2115_;
  assign po084 = new_n1300_ | new_n1312_;
  assign new_n1314_ = new_n1481_ & pi141 & new_n2115_;
  assign po085 = new_n1301_ | new_n1314_;
  assign new_n1316_ = new_n1481_ & pi142 & new_n2115_;
  assign po086 = new_n1302_ | new_n1316_;
  assign new_n1318_ = new_n1481_ & pi143 & new_n2115_;
  assign po087 = new_n1303_ | new_n1318_;
  assign new_n1320_ = new_n1481_ & pi144 & new_n2115_;
  assign po088 = new_n1304_ | new_n1320_;
  assign new_n1322_ = new_n1481_ & pi145 & new_n2115_;
  assign po089 = new_n1305_ | new_n1322_;
  assign new_n1324_ = new_n1481_ & pi146 & new_n2115_;
  assign po090 = new_n1306_ | new_n1324_;
  assign new_n1326_ = new_n1481_ & pi147 & new_n2115_;
  assign po091 = new_n1307_ | new_n1326_;
  assign new_n1328_ = new_n2116_ & new_n1486_ & new_n1210_ & new_n2097_ & new_n2098_ & new_n1102_ & new_n2108_ & new_n1485_;
  assign new_n1329_ = new_n2116_ & new_n1486_ & new_n1210_ & new_n2097_ & new_n2098_ & new_n1104_ & new_n2108_ & new_n1485_;
  assign new_n1330_ = new_n2116_ & new_n1486_ & new_n1210_ & new_n2097_ & new_n2098_ & new_n1106_ & new_n2108_ & new_n1485_;
  assign new_n1331_ = new_n2116_ & new_n1486_ & new_n1210_ & new_n2097_ & new_n2098_ & new_n1108_ & new_n2108_ & new_n1485_;
  assign new_n1332_ = new_n1481_ & pi003 & new_n2117_;
  assign new_n1333_ = new_n1328_ | new_n1332_;
  assign new_n1334_ = new_n1481_ & pi002 & new_n2117_;
  assign new_n1335_ = new_n1329_ | new_n1334_;
  assign new_n1336_ = new_n1481_ & pi001 & new_n2117_;
  assign new_n1337_ = new_n1330_ | new_n1336_;
  assign new_n1338_ = new_n1481_ & pi000 & new_n2117_;
  assign new_n1339_ = new_n1331_ | new_n1338_;
  assign po092 = pi148 & new_n530_;
  assign po093 = new_n1627_ & new_n1625_ & new_n1623_ & new_n1624_ & new_n1626_ & pi148 & pi072;
  assign po094 = pi148 & pi052;
  assign po095 = pi149 & pi052;
  assign po096 = pi149 & pi073;
  assign po097 = new_n1359_ & po096;
  assign po098 = pi074 & new_n530_;
  assign po099 = pi074 & pi052;
  assign po100 = pi074 & pi072;
  assign po101 = pi069 & po100;
  assign po102 = pi074 & pi073;
  assign po103 = pi148 & pi073;
  assign new_n1352_ = new_n902_ | new_n644_ | new_n861_ | new_n860_ | new_n854_ | new_n558_ | new_n859_;
  assign new_n1353_ = ~new_n1352_;
  assign new_n1354_ = ~new_n900_;
  assign new_n1355_ = ~new_n901_;
  assign new_n1356_ = pi014 & new_n645_ & new_n641_ & new_n1049_;
  assign new_n1357_ = new_n641_ & new_n1049_ & new_n887_ & new_n1354_ & new_n1353_ & new_n1355_ & new_n1754_ & pi015;
  assign po104 = new_n1356_ | new_n1357_;
  assign new_n1359_ = ~pi014;
  assign new_n1360_ = new_n868_ & pi004;
  assign new_n1361_ = ~new_n1360_;
  assign new_n1362_ = ~new_n1982_;
  assign new_n1363_ = new_n2118_ & new_n1362_ & pi151 & new_n1361_ & pi150;
  assign new_n1364_ = new_n1982_ & new_n1610_ & new_n2119_;
  assign po105 = new_n1363_ | new_n1364_;
  assign new_n1366_ = ~new_n1977_;
  assign new_n1367_ = new_n2120_ & new_n1366_ & pi152 & new_n1361_ & pi150;
  assign new_n1368_ = new_n2120_ & new_n1366_ & pi153 & new_n1361_ & pi150;
  assign new_n1369_ = new_n2120_ & new_n1366_ & pi154 & new_n1361_ & pi150;
  assign new_n1370_ = new_n2120_ & new_n1366_ & pi155 & new_n1361_ & pi150;
  assign new_n1371_ = new_n2120_ & new_n1366_ & pi156 & new_n1361_ & pi150;
  assign new_n1372_ = new_n1977_ & pi063 & new_n2121_;
  assign po106 = new_n1367_ | new_n1372_;
  assign new_n1374_ = new_n1977_ & pi062 & new_n2121_;
  assign po107 = new_n1368_ | new_n1374_;
  assign new_n1376_ = new_n1977_ & pi061 & new_n2121_;
  assign po108 = new_n1369_ | new_n1376_;
  assign new_n1378_ = new_n1977_ & pi060 & new_n2121_;
  assign po109 = new_n1370_ | new_n1378_;
  assign new_n1380_ = new_n1977_ & pi075 & new_n2121_;
  assign po110 = new_n1371_ | new_n1380_;
  assign new_n1382_ = new_n1855_ & new_n2908_;
  assign new_n1383_ = new_n1857_ & new_n1382_;
  assign new_n1384_ = new_n2923_ & new_n1382_;
  assign new_n1385_ = new_n2923_ & new_n1857_;
  assign new_n1386_ = new_n1384_ | new_n1385_ | new_n1383_;
  assign new_n1387_ = new_n1848_ & new_n1386_;
  assign new_n1388_ = new_n2928_ & new_n1386_;
  assign new_n1389_ = new_n2928_ & new_n1848_;
  assign new_n1390_ = new_n1388_ | new_n1389_ | new_n1387_;
  assign new_n1391_ = ~new_n2598_;
  assign new_n1392_ = ~new_n2613_;
  assign new_n1393_ = ~new_n2618_;
  assign new_n1394_ = new_n1392_ & new_n1391_;
  assign new_n1395_ = new_n1393_ & new_n1394_;
  assign new_n1396_ = ~new_n1391_;
  assign new_n1397_ = ~new_n2628_;
  assign new_n1398_ = ~new_n2633_;
  assign new_n1399_ = new_n1397_ & new_n1396_;
  assign new_n1400_ = new_n1398_ & new_n1399_;
  assign new_n1401_ = new_n2122_ & new_n2623_ & new_n1857_;
  assign new_n1402_ = new_n1869_ & new_n2653_ & new_n2123_;
  assign new_n1403_ = new_n1401_ | new_n1402_;
  assign new_n1404_ = new_n2124_ & new_n2618_ & new_n1857_;
  assign new_n1405_ = new_n1869_ & new_n2648_ & new_n2125_;
  assign new_n1406_ = new_n1404_ | new_n1405_;
  assign new_n1407_ = new_n2126_ & new_n2613_ & new_n1857_;
  assign new_n1408_ = new_n1869_ & new_n2643_ & new_n2127_;
  assign new_n1409_ = new_n1407_ | new_n1408_;
  assign new_n1410_ = new_n2128_ & new_n2598_ & new_n1857_;
  assign new_n1411_ = new_n1869_ & new_n1396_ & new_n2129_;
  assign new_n1412_ = new_n1410_ | new_n1411_;
  assign new_n1413_ = ~new_n1412_;
  assign new_n1414_ = ~new_n1409_;
  assign new_n1415_ = ~new_n1406_;
  assign new_n1416_ = new_n1414_ & new_n1413_;
  assign new_n1417_ = new_n1415_ & new_n1416_;
  assign new_n1418_ = new_n2130_ & new_n2623_ & new_n1855_;
  assign new_n1419_ = new_n1868_ & new_n2668_ & new_n2131_;
  assign new_n1420_ = new_n1418_ | new_n1419_;
  assign new_n1421_ = new_n2132_ & new_n2618_ & new_n1855_;
  assign new_n1422_ = new_n1868_ & new_n2663_ & new_n2133_;
  assign new_n1423_ = new_n1421_ | new_n1422_;
  assign new_n1424_ = new_n2134_ & new_n2613_ & new_n1855_;
  assign new_n1425_ = new_n1868_ & new_n2658_ & new_n2135_;
  assign new_n1426_ = new_n1424_ | new_n1425_;
  assign new_n1427_ = new_n2136_ & new_n2598_ & new_n1855_;
  assign new_n1428_ = new_n1868_ & new_n1413_ & new_n2137_;
  assign new_n1429_ = new_n1427_ | new_n1428_;
  assign new_n1430_ = ~new_n867_;
  assign new_n1431_ = ~new_n657_;
  assign new_n1432_ = ~new_n864_;
  assign new_n1433_ = ~new_n871_;
  assign po111 = pi014 & new_n937_ & new_n1432_ & new_n1430_ & new_n926_ & new_n1431_ & new_n1433_ & new_n938_ & new_n641_ & new_n1049_;
  assign new_n1435_ = pi161 & pi160 & pi159 & pi157 & pi158;
  assign new_n1436_ = pi161 & pi160 & pi157 & pi158;
  assign new_n1437_ = pi161 & pi157 & pi158;
  assign new_n1438_ = pi157 & pi161;
  assign po112 = ~pi157;
  assign new_n1440_ = ~new_n2006_;
  assign new_n1441_ = ~new_n532_;
  assign po113 = new_n1440_ & new_n1441_ & new_n918_;
  assign new_n1443_ = ~new_n2016_;
  assign po114 = new_n1443_ & new_n1441_ & new_n918_;
  assign new_n1445_ = ~new_n539_;
  assign po115 = new_n1441_ & new_n1445_ & new_n918_;
  assign new_n1447_ = ~new_n500_;
  assign po116 = new_n1441_ & new_n1447_ & new_n918_;
  assign new_n1449_ = ~new_n1846_;
  assign po117 = new_n1441_ & new_n1449_ & new_n918_;
  assign po118 = pi052 & pi162;
  assign new_n1452_ = ~new_n559_;
  assign new_n1453_ = ~new_n874_;
  assign new_n1454_ = new_n1452_ & pi077 & new_n1453_ & new_n641_ & new_n1049_;
  assign new_n1455_ = pi019 & pi062 & new_n824_ & pi075 & new_n825_ & po052 & new_n641_ & new_n1049_;
  assign po119 = new_n1455_ | new_n1454_;
  assign new_n1457_ = new_n902_ & new_n1510_;
  assign new_n1458_ = pi163 | pi015 | pi004;
  assign new_n1459_ = new_n834_ | new_n833_;
  assign new_n1460_ = pi015 | pi163;
  assign new_n1461_ = new_n862_ | new_n854_ | new_n843_ | new_n1457_ | new_n864_;
  assign new_n1462_ = pi165 | pi004 | pi164;
  assign new_n1463_ = new_n902_ | new_n854_;
  assign new_n1464_ = ~new_n860_;
  assign new_n1465_ = ~new_n859_;
  assign new_n1466_ = po052 & new_n1458_;
  assign new_n1467_ = new_n860_ & new_n1509_;
  assign new_n1468_ = new_n1460_ & new_n860_ & new_n1510_;
  assign new_n1469_ = ~new_n1479_;
  assign new_n1470_ = new_n1462_ & new_n1469_ & new_n1461_;
  assign new_n1471_ = pi163 & new_n1463_;
  assign new_n1472_ = ~new_n1466_;
  assign new_n1473_ = new_n859_ | new_n902_ | new_n1459_;
  assign new_n1474_ = ~new_n1471_;
  assign new_n1475_ = pi004 & new_n645_;
  assign new_n1476_ = pi163 & new_n645_;
  assign new_n1477_ = pi004 & new_n569_;
  assign new_n1478_ = pi163 & new_n569_;
  assign new_n1479_ = new_n1475_ | new_n1477_ | new_n1478_ | new_n1476_;
  assign new_n1480_ = new_n1052_ & pi164 & new_n1464_ & new_n926_ & new_n1465_;
  assign new_n1481_ = new_n1480_ | new_n878_ | new_n1470_;
  assign new_n1482_ = new_n898_ & new_n1473_;
  assign new_n1483_ = ~new_n1481_;
  assign new_n1484_ = ~new_n1474_;
  assign new_n1485_ = new_n1468_ | new_n1482_ | new_n1467_;
  assign new_n1486_ = new_n1484_ | new_n1483_;
  assign po120 = pi030 & pi052;
  assign new_n1488_ = ~new_n723_;
  assign new_n1489_ = new_n919_ & new_n1488_;
  assign po121 = new_n1488_ & new_n1441_;
  assign new_n1491_ = new_n791_ & pi166;
  assign po122 = pi073 & pi030;
  assign po123 = pi072 & pi030;
  assign new_n1494_ = ~new_n1491_;
  assign po124 = new_n1494_ & new_n919_ & new_n1488_;
  assign po125 = new_n641_ & pi018 & new_n1049_;
  assign new_n1497_ = ~new_n902_;
  assign new_n1498_ = ~new_n1505_;
  assign new_n1499_ = new_n641_ & new_n1498_ & new_n1497_;
  assign new_n1500_ = pi167 & new_n902_;
  assign new_n1501_ = new_n1506_ | new_n1500_;
  assign new_n1502_ = pi150 & new_n1501_;
  assign po126 = new_n879_ | new_n1499_;
  assign po127 = ~new_n1502_;
  assign new_n1505_ = ~pi167;
  assign new_n1506_ = ~pi168;
  assign new_n1507_ = new_n902_ & pi167;
  assign new_n1508_ = ~new_n1507_;
  assign new_n1509_ = pi168 & new_n1508_;
  assign new_n1510_ = ~new_n1509_;
  assign new_n1511_ = new_n1845_ | new_n1839_;
  assign new_n1512_ = new_n1516_ & new_n1511_ & pi150;
  assign new_n1513_ = ~new_n1511_;
  assign new_n1514_ = pi084 & new_n1513_ & pi150;
  assign po128 = new_n1514_ | new_n1512_;
  assign new_n1516_ = ~pi084;
  assign new_n1517_ = new_n1839_ & pi084;
  assign new_n1518_ = new_n1845_ & new_n1516_;
  assign new_n1519_ = new_n1518_ | new_n1517_;
  assign new_n1520_ = pi150 & new_n1524_ & new_n1519_;
  assign new_n1521_ = ~new_n1519_;
  assign new_n1522_ = pi150 & pi169 & new_n1521_;
  assign po129 = new_n1522_ | new_n1520_;
  assign new_n1524_ = ~pi169;
  assign new_n1525_ = new_n1517_ & pi169;
  assign new_n1526_ = new_n1518_ & new_n1524_;
  assign new_n1527_ = new_n1526_ | new_n1525_;
  assign new_n1528_ = pi150 & new_n1532_ & new_n1527_;
  assign new_n1529_ = ~new_n1527_;
  assign new_n1530_ = pi150 & pi170 & new_n1529_;
  assign po130 = new_n1530_ | new_n1528_;
  assign new_n1532_ = ~pi170;
  assign new_n1533_ = ~new_n870_;
  assign po131 = pi171 & new_n1049_ & new_n1533_ & new_n641_;
  assign new_n1535_ = new_n902_ | new_n834_ | new_n899_;
  assign new_n1536_ = new_n877_ | new_n872_ | new_n878_;
  assign new_n1537_ = po065 & new_n1535_;
  assign new_n1538_ = pi004 & new_n1536_;
  assign new_n1539_ = new_n1538_ | new_n1537_;
  assign new_n1540_ = new_n1645_ & new_n1539_;
  assign new_n1541_ = ~new_n834_;
  assign new_n1542_ = new_n1541_ & po165;
  assign new_n1543_ = new_n834_ & po065 & po165;
  assign po132 = new_n1542_ | new_n1543_ | new_n1540_;
  assign po133 = ~pi021;
  assign new_n1546_ = ~pi018;
  assign new_n1547_ = ~pi172;
  assign new_n1548_ = ~pi173;
  assign new_n1549_ = ~pi019;
  assign new_n1550_ = new_n1548_ & new_n1546_ & new_n1549_ & new_n1547_;
  assign new_n1551_ = ~new_n1550_;
  assign new_n1552_ = ~new_n1995_;
  assign new_n1553_ = ~new_n1557_;
  assign new_n1554_ = new_n1552_ & new_n1551_ & new_n1553_ & new_n641_;
  assign new_n1555_ = pi017 & pi018;
  assign po134 = new_n1558_ | new_n1554_;
  assign new_n1557_ = ~pi017;
  assign new_n1558_ = po133 & pi174;
  assign po135 = ~pi175;
  assign new_n1560_ = ~new_n1998_;
  assign new_n1561_ = new_n676_ & new_n504_ & new_n1560_;
  assign new_n1562_ = ~new_n1561_;
  assign new_n1563_ = ~new_n1998_;
  assign new_n1564_ = ~new_n504_;
  assign new_n1565_ = new_n1564_ & new_n1563_;
  assign new_n1566_ = ~new_n1565_;
  assign new_n1567_ = po139 & new_n1560_;
  assign new_n1568_ = po139 & new_n1562_;
  assign new_n1569_ = po139 & new_n1566_;
  assign new_n1570_ = ~po139;
  assign new_n1571_ = new_n1570_ & new_n529_;
  assign po136 = new_n1567_ | new_n1571_;
  assign new_n1573_ = new_n1570_ & new_n528_;
  assign po137 = new_n1568_ | new_n1573_;
  assign new_n1575_ = new_n1570_ & new_n527_;
  assign po138 = new_n1569_ | new_n1575_;
  assign new_n1577_ = new_n2007_ & pi168;
  assign new_n1578_ = ~pi176;
  assign new_n1579_ = ~pi042;
  assign new_n1580_ = new_n1579_ & new_n640_;
  assign new_n1581_ = pi004 & pi177;
  assign new_n1582_ = pi178 & pi004 & new_n1459_;
  assign new_n1583_ = ~new_n1578_;
  assign new_n1584_ = ~pi012;
  assign new_n1585_ = ~new_n1577_;
  assign new_n1586_ = ~new_n1581_;
  assign new_n1587_ = ~new_n1582_;
  assign new_n1588_ = new_n1586_ & new_n1584_ & new_n1583_ & new_n1587_ & new_n1585_;
  assign new_n1589_ = ~pi177;
  assign new_n1590_ = new_n1589_ & new_n564_;
  assign new_n1591_ = pi015 & new_n657_;
  assign new_n1592_ = ~new_n1580_;
  assign new_n1593_ = ~new_n1588_;
  assign new_n1594_ = ~new_n1590_;
  assign new_n1595_ = ~new_n1591_;
  assign new_n1596_ = new_n1594_ & new_n1592_ & new_n1595_ & new_n1593_;
  assign new_n1597_ = ~new_n1596_;
  assign new_n1598_ = ~new_n676_;
  assign new_n1599_ = new_n1598_ & new_n1563_ & new_n1597_;
  assign po139 = ~new_n1599_;
  assign po140 = new_n641_ & pi172 & new_n1049_;
  assign new_n1602_ = pi179 | pi173;
  assign po141 = new_n641_ & new_n1602_ & new_n1049_;
  assign new_n1604_ = ~pi075;
  assign new_n1605_ = ~pi060;
  assign new_n1606_ = ~pi061;
  assign new_n1607_ = ~pi062;
  assign new_n1608_ = ~pi063;
  assign new_n1609_ = new_n1607_ & new_n1605_ & new_n1604_ & new_n1608_ & new_n1606_;
  assign new_n1610_ = new_n1680_ | new_n1609_;
  assign new_n1611_ = new_n2138_ & new_n854_ & new_n1983_ & new_n936_;
  assign new_n1612_ = new_n2138_ & new_n854_ & new_n2898_ & new_n936_;
  assign new_n1613_ = new_n537_ & po082 & new_n2139_;
  assign po142 = new_n1611_ | new_n1613_;
  assign new_n1615_ = new_n537_ & po083 & new_n2139_;
  assign po143 = new_n1612_ | new_n1615_;
  assign new_n1617_ = pi180 | pi163;
  assign new_n1618_ = new_n902_ | new_n843_ | new_n864_ | new_n862_ | new_n863_ | new_n854_;
  assign new_n1619_ = pi165 & new_n1618_;
  assign new_n1620_ = ~pi165;
  assign new_n1621_ = new_n1620_ & new_n872_;
  assign new_n1622_ = new_n1617_ & new_n878_;
  assign new_n1623_ = ~new_n1619_;
  assign new_n1624_ = ~new_n1621_;
  assign new_n1625_ = ~new_n1622_;
  assign new_n1626_ = ~pi016;
  assign new_n1627_ = ~pi008;
  assign new_n1628_ = pi043 & pi181;
  assign new_n1629_ = ~new_n1628_;
  assign new_n1630_ = ~po186;
  assign new_n1631_ = ~new_n1754_;
  assign new_n1632_ = new_n1631_ & new_n1630_;
  assign new_n1633_ = po160 & new_n830_;
  assign new_n1634_ = new_n831_ & po160;
  assign new_n1635_ = po160 & new_n552_ & new_n1876_;
  assign new_n1636_ = pi037 & po160 & new_n552_ & new_n745_;
  assign new_n1637_ = ~new_n1635_;
  assign new_n1638_ = ~new_n550_;
  assign new_n1639_ = ~new_n1632_;
  assign new_n1640_ = ~new_n1633_;
  assign new_n1641_ = ~new_n1634_;
  assign new_n1642_ = ~new_n1636_;
  assign new_n1643_ = ~new_n2768_;
  assign new_n1644_ = ~new_n2773_;
  assign new_n1645_ = new_n1644_ | new_n1643_;
  assign po144 = ~new_n2838_;
  assign po145 = ~new_n2843_;
  assign new_n1648_ = pi182 & po186;
  assign new_n1649_ = new_n828_ & pi016;
  assign new_n1650_ = new_n1998_ & pi016;
  assign new_n1651_ = ~new_n932_;
  assign new_n1652_ = ~pi183;
  assign new_n1653_ = ~pi182;
  assign po146 = new_n1648_ | new_n1650_ | new_n932_ | new_n1649_;
  assign new_n1655_ = pi015 & pi184;
  assign new_n1656_ = pi014 & pi185;
  assign new_n1657_ = new_n1656_ | new_n1655_;
  assign new_n1658_ = new_n872_ & new_n1657_;
  assign new_n1659_ = ~pi186;
  assign new_n1660_ = ~new_n751_;
  assign new_n1661_ = ~new_n874_;
  assign new_n1662_ = new_n1660_ & new_n1661_ & new_n1659_;
  assign po147 = new_n1662_ | new_n762_ | new_n1658_;
  assign new_n1664_ = ~pi150;
  assign new_n1665_ = new_n902_ | new_n899_;
  assign new_n1666_ = new_n874_ | new_n872_ | new_n901_ | new_n873_;
  assign new_n1667_ = new_n897_ & po065 & new_n1665_;
  assign new_n1668_ = new_n834_ & po065;
  assign new_n1669_ = pi018 & new_n870_;
  assign new_n1670_ = pi004 & new_n1666_;
  assign new_n1671_ = po052 & pi018;
  assign new_n1672_ = pi026 & po065 & new_n834_;
  assign new_n1673_ = new_n820_ & new_n899_;
  assign new_n1674_ = po186 & new_n834_;
  assign new_n1675_ = new_n1668_ | new_n1670_ | new_n1667_ | new_n1671_ | new_n1669_;
  assign new_n1676_ = new_n1673_ | new_n871_ | new_n1674_ | new_n901_;
  assign new_n1677_ = new_n494_ & new_n1675_;
  assign new_n1678_ = new_n496_ & new_n1680_ & new_n1676_ & pi150 & new_n502_;
  assign po148 = new_n1677_ | new_n1672_ | new_n1678_;
  assign new_n1680_ = pi187 & new_n1586_;
  assign new_n1681_ = new_n860_ | new_n859_ | new_n902_;
  assign new_n1682_ = new_n1509_ & new_n1681_;
  assign new_n1683_ = ~new_n1682_;
  assign new_n1684_ = ~pi078;
  assign new_n1685_ = new_n1684_ & pi188 & new_n1683_ & new_n557_ & new_n502_ & new_n1719_;
  assign po149 = ~new_n1685_;
  assign new_n1687_ = new_n875_ | new_n868_ | new_n1721_ | new_n877_ | new_n879_ | new_n869_ | new_n876_;
  assign new_n1688_ = ~new_n1687_;
  assign new_n1689_ = ~new_n1721_;
  assign new_n1690_ = new_n1661_ & new_n1689_ & new_n1688_ & new_n938_ & new_n937_;
  assign new_n1691_ = ~new_n1690_;
  assign new_n1692_ = ~new_n945_;
  assign new_n1693_ = ~new_n829_;
  assign new_n1694_ = new_n1693_ & new_n1691_ & new_n1563_ & new_n502_ & new_n1692_;
  assign new_n1695_ = ~new_n1780_;
  assign new_n1696_ = new_n1695_ & new_n502_ & new_n1688_;
  assign new_n1697_ = new_n936_ & new_n502_ & new_n831_;
  assign new_n1698_ = new_n870_ & pi018;
  assign new_n1699_ = ~new_n1694_;
  assign new_n1700_ = ~new_n1696_;
  assign new_n1701_ = ~new_n1697_;
  assign new_n1702_ = ~new_n1698_;
  assign po150 = new_n1701_ & new_n1699_ & new_n1702_ & new_n1700_;
  assign new_n1704_ = ~pi189;
  assign po151 = ~pi190;
  assign new_n1706_ = pi059 & pi064 & pi058 & new_n1704_ & pi191 & pi060 & pi075 & pi061 & pi063 & pi062;
  assign new_n1707_ = po052 & pi059 & pi064 & pi058 & pi062 & pi060 & pi075 & pi061 & pi191 & pi019 & pi063;
  assign new_n1708_ = new_n1707_ | new_n1706_;
  assign new_n1709_ = pi084 & new_n1532_ & new_n1072_ & new_n1524_;
  assign new_n1710_ = ~new_n1714_;
  assign new_n1711_ = ~new_n1709_;
  assign new_n1712_ = new_n1711_ & new_n641_ & new_n1710_;
  assign po152 = new_n1712_ | new_n1708_;
  assign new_n1714_ = ~pi192;
  assign new_n1715_ = new_n1708_ | pi192;
  assign new_n1716_ = ~new_n1712_;
  assign new_n1717_ = new_n1844_ & new_n1710_ & new_n1716_;
  assign new_n1718_ = ~new_n1717_;
  assign new_n1719_ = ~new_n1715_;
  assign new_n1720_ = new_n1712_ & pi192;
  assign new_n1721_ = new_n1708_ | new_n1720_;
  assign new_n1722_ = new_n869_ & pi004;
  assign new_n1723_ = ~new_n1722_;
  assign new_n1724_ = ~new_n1981_;
  assign new_n1725_ = new_n2140_ & new_n1724_ & pi193 & new_n1723_ & pi150;
  assign new_n1726_ = new_n1981_ & new_n1610_ & new_n2141_;
  assign po153 = new_n1725_ | new_n1726_;
  assign new_n1728_ = ~new_n1976_;
  assign new_n1729_ = new_n2142_ & new_n1728_ & pi194 & new_n1723_ & pi150;
  assign new_n1730_ = new_n2142_ & new_n1728_ & pi195 & new_n1723_ & pi150;
  assign new_n1731_ = new_n2142_ & new_n1728_ & pi196 & new_n1723_ & pi150;
  assign new_n1732_ = new_n2142_ & new_n1728_ & pi197 & new_n1723_ & pi150;
  assign new_n1733_ = new_n2142_ & new_n1728_ & pi198 & new_n1723_ & pi150;
  assign new_n1734_ = new_n1976_ & pi063 & new_n2143_;
  assign po154 = new_n1729_ | new_n1734_;
  assign new_n1736_ = new_n1976_ & pi062 & new_n2143_;
  assign po155 = new_n1730_ | new_n1736_;
  assign new_n1738_ = new_n1976_ & pi061 & new_n2143_;
  assign po156 = new_n1731_ | new_n1738_;
  assign new_n1740_ = new_n1976_ & pi060 & new_n2143_;
  assign po157 = new_n1732_ | new_n1740_;
  assign new_n1742_ = new_n1976_ & pi075 & new_n2143_;
  assign po158 = new_n1733_ | new_n1742_;
  assign new_n1744_ = new_n960_ & new_n854_;
  assign new_n1745_ = new_n854_ | new_n579_;
  assign new_n1746_ = po065 & new_n1745_;
  assign new_n1747_ = ~new_n1744_;
  assign new_n1748_ = ~new_n1752_;
  assign new_n1749_ = ~new_n830_;
  assign new_n1750_ = new_n1589_ & new_n1748_ & new_n1747_ & new_n1049_ & new_n496_ & new_n1749_;
  assign po159 = new_n1750_ | new_n1746_;
  assign new_n1752_ = ~pi199;
  assign po160 = new_n1589_ & new_n496_ & pi199;
  assign new_n1754_ = ~po160;
  assign new_n1755_ = pi128 & new_n1876_;
  assign new_n1756_ = ~po139;
  assign new_n1757_ = new_n1756_ & new_n2007_ & new_n1755_;
  assign new_n1758_ = ~new_n2003_;
  assign new_n1759_ = new_n1758_ & new_n641_ & pi200;
  assign po161 = new_n1759_ | new_n1757_;
  assign new_n1761_ = ~new_n1755_;
  assign new_n1762_ = new_n860_ | new_n902_;
  assign new_n1763_ = pi201 & new_n1762_;
  assign new_n1764_ = new_n866_ & new_n1433_ & new_n1355_ & new_n1541_ & new_n1680_;
  assign new_n1765_ = pi015 & new_n1680_ & new_n1541_ & new_n820_;
  assign new_n1766_ = new_n901_ & new_n1680_ & new_n1541_ & pi015;
  assign new_n1767_ = pi014 & new_n1680_ & new_n1541_ & new_n871_;
  assign new_n1768_ = ~new_n1763_;
  assign new_n1769_ = new_n1465_ & new_n1768_;
  assign po162 = new_n1781_ & new_n936_ & new_n1769_ & new_n502_ & new_n831_;
  assign new_n1771_ = ~new_n1769_;
  assign new_n1772_ = new_n496_ & new_n1764_;
  assign new_n1773_ = new_n496_ & new_n1765_;
  assign new_n1774_ = new_n1766_ & new_n496_;
  assign po163 = new_n1772_ | new_n1774_ | new_n1782_ | new_n1767_ | new_n1773_;
  assign new_n1776_ = ~new_n858_;
  assign new_n1777_ = ~new_n880_;
  assign new_n1778_ = new_n1776_ & pi005 & new_n1777_ & pi202;
  assign po164 = ~new_n1778_;
  assign new_n1780_ = ~po163;
  assign new_n1781_ = ~pi078;
  assign new_n1782_ = new_n828_ & pi078;
  assign new_n1783_ = pi004 & new_n884_;
  assign new_n1784_ = pi203 & pi204;
  assign new_n1785_ = new_n1875_ & pi204;
  assign new_n1786_ = pi203 & new_n1874_;
  assign new_n1787_ = ~new_n1783_;
  assign new_n1788_ = new_n833_ & new_n1786_;
  assign new_n1789_ = pi150 & pi205 & new_n1787_;
  assign new_n1790_ = new_n858_ & new_n1786_;
  assign po165 = new_n1785_ | new_n1784_;
  assign po166 = new_n1786_ | new_n1785_;
  assign po167 = new_n1789_ | new_n1790_ | new_n1788_;
  assign po168 = ~pi205;
  assign new_n1795_ = ~new_n878_;
  assign new_n1796_ = new_n2144_ & new_n2146_ & new_n878_;
  assign new_n1797_ = new_n2144_ & new_n2145_ & new_n878_;
  assign new_n1798_ = new_n1795_ & new_n2149_ & new_n2147_;
  assign po169 = new_n1796_ | new_n1798_;
  assign new_n1800_ = new_n1795_ & new_n2148_ & new_n2147_;
  assign po170 = new_n1797_ | new_n1800_;
  assign new_n1802_ = new_n2150_ & new_n2152_ & new_n1795_;
  assign new_n1803_ = new_n2150_ & new_n2151_ & new_n1795_;
  assign new_n1804_ = new_n878_ & new_n2155_ & new_n2153_;
  assign po171 = new_n1802_ | new_n1804_;
  assign new_n1806_ = new_n878_ & new_n2154_ & new_n2153_;
  assign po172 = new_n1803_ | new_n1806_;
  assign new_n1808_ = ~po079;
  assign new_n1809_ = new_n2156_ & new_n2165_ & pi022;
  assign new_n1810_ = new_n2156_ & new_n2164_ & pi022;
  assign new_n1811_ = new_n2156_ & new_n2163_ & pi022;
  assign new_n1812_ = new_n2156_ & new_n2162_ & pi022;
  assign new_n1813_ = new_n2156_ & new_n2161_ & pi022;
  assign new_n1814_ = new_n2156_ & new_n2160_ & pi022;
  assign new_n1815_ = new_n2156_ & new_n2159_ & pi022;
  assign new_n1816_ = new_n2156_ & new_n2158_ & pi022;
  assign new_n1817_ = new_n2156_ & new_n2157_ & pi022;
  assign new_n1818_ = new_n2156_ & new_n1808_ & pi022;
  assign new_n1819_ = new_n594_ & po000 & new_n2166_;
  assign po173 = new_n1809_ | new_n1819_;
  assign new_n1821_ = new_n594_ & new_n2174_ & new_n2166_;
  assign po174 = new_n1810_ | new_n1821_;
  assign new_n1823_ = new_n594_ & new_n2173_ & new_n2166_;
  assign po175 = new_n1811_ | new_n1823_;
  assign new_n1825_ = new_n594_ & new_n2172_ & new_n2166_;
  assign po176 = new_n1812_ | new_n1825_;
  assign new_n1827_ = new_n594_ & new_n2171_ & new_n2166_;
  assign po177 = new_n1813_ | new_n1827_;
  assign new_n1829_ = new_n594_ & new_n2170_ & new_n2166_;
  assign po178 = new_n1814_ | new_n1829_;
  assign new_n1831_ = new_n594_ & new_n2169_ & new_n2166_;
  assign po179 = new_n1815_ | new_n1831_;
  assign new_n1833_ = new_n594_ & new_n2168_ & new_n2166_;
  assign po180 = new_n1816_ | new_n1833_;
  assign new_n1835_ = new_n594_ & new_n2167_ & new_n2166_;
  assign po181 = new_n1817_ | new_n1835_;
  assign new_n1837_ = new_n594_ & po000 & new_n2166_;
  assign po182 = new_n1818_ | new_n1837_;
  assign new_n1839_ = pi206 & new_n1435_;
  assign new_n1840_ = new_n1843_ | new_n1839_;
  assign po183 = pi150 & new_n1840_;
  assign po184 = ~pi191;
  assign new_n1843_ = new_n1718_ & pi191;
  assign new_n1844_ = pi014 | pi179 | pi004;
  assign new_n1845_ = new_n1715_ & new_n1844_;
  assign new_n1846_ = ~new_n1845_;
  assign new_n1847_ = pi207 & pi083;
  assign new_n1848_ = pi208 & pi082;
  assign new_n1849_ = pi209 & pi081;
  assign new_n1850_ = ~pi081;
  assign new_n1851_ = pi209 & new_n1850_;
  assign new_n1852_ = ~pi209;
  assign new_n1853_ = new_n1852_ & pi081;
  assign new_n1854_ = ~pi082;
  assign new_n1855_ = pi208 & new_n1854_;
  assign new_n1856_ = ~pi208;
  assign new_n1857_ = new_n1856_ & pi082;
  assign new_n1858_ = ~pi083;
  assign new_n1859_ = pi207 & new_n1858_;
  assign new_n1860_ = ~pi207;
  assign new_n1861_ = new_n1860_ & pi083;
  assign new_n1862_ = pi207 | pi083;
  assign new_n1863_ = pi208 | pi082;
  assign new_n1864_ = pi209 | pi081;
  assign new_n1865_ = pi011 | pi010;
  assign new_n1866_ = ~new_n1851_;
  assign new_n1867_ = ~new_n1853_;
  assign new_n1868_ = ~new_n1855_;
  assign new_n1869_ = ~new_n1857_;
  assign new_n1870_ = ~new_n1859_;
  assign new_n1871_ = ~new_n1861_;
  assign po185 = ~pi210;
  assign po186 = ~pi039;
  assign new_n1874_ = ~pi204;
  assign new_n1875_ = ~pi203;
  assign new_n1876_ = pi120 & pi122 & pi124 & pi126 & pi127 & pi125 & pi123 & pi119 & pi121;
  assign new_n1877_ = pi120 & pi122 & pi124 & pi126 & pi125 & pi123 & pi119 & pi121;
  assign new_n1878_ = pi120 & pi122 & pi124 & pi125 & pi123 & pi119 & pi121;
  assign new_n1879_ = pi120 & pi122 & pi124 & pi123 & pi119 & pi121;
  assign new_n1880_ = pi120 & pi122 & pi123 & pi119 & pi121;
  assign new_n1881_ = pi120 & pi122 & pi119 & pi121;
  assign new_n1882_ = pi120 & pi119 & pi121;
  assign new_n1883_ = pi119 & pi120;
  assign new_n1884_ = ~pi119;
  assign new_n1885_ = new_n902_ & new_n1540_;
  assign new_n1886_ = new_n858_ & new_n1991_;
  assign new_n1887_ = new_n833_ & new_n1991_;
  assign new_n1888_ = ~new_n1902_;
  assign new_n1889_ = pi211 & new_n1888_;
  assign new_n1890_ = pi212 & new_n1888_;
  assign new_n1891_ = pi213 & new_n1888_;
  assign new_n1892_ = pi214 & new_n1888_;
  assign new_n1893_ = pi215 & new_n1888_;
  assign new_n1894_ = ~new_n1783_;
  assign new_n1895_ = pi216 & new_n1894_;
  assign po187 = new_n1784_ | new_n1889_ | new_n1540_;
  assign po188 = new_n1885_ | new_n1890_;
  assign po189 = new_n1886_ | new_n1891_;
  assign po190 = new_n1887_ | new_n1892_;
  assign po191 = new_n1785_ | new_n1893_;
  assign po192 = new_n1786_ | new_n1895_;
  assign new_n1902_ = pi004 & new_n883_;
  assign new_n1903_ = new_n2176_ & new_n2177_ & new_n2178_ & pi194 & new_n869_;
  assign new_n1904_ = new_n2176_ & new_n2177_ & new_n2178_ & pi195 & new_n869_;
  assign new_n1905_ = new_n2176_ & new_n2177_ & new_n2178_ & pi196 & new_n869_;
  assign new_n1906_ = new_n2176_ & new_n2177_ & new_n2178_ & pi197 & new_n869_;
  assign new_n1907_ = new_n2176_ & new_n2177_ & new_n2178_ & pi198 & new_n869_;
  assign new_n1908_ = new_n2176_ & new_n2177_ & new_n2178_ & pi193 & new_n869_;
  assign new_n1909_ = new_n2179_ & new_n2180_ & new_n868_ & pi152 & new_n2181_;
  assign po193 = new_n1921_ | new_n1903_ | new_n1909_;
  assign new_n1911_ = new_n2179_ & new_n2180_ & new_n868_ & pi153 & new_n2181_;
  assign po194 = new_n1922_ | new_n1927_ | new_n1904_ | new_n1911_;
  assign new_n1913_ = new_n2179_ & new_n2180_ & new_n868_ & pi154 & new_n2181_;
  assign po195 = new_n1923_ | new_n1928_ | new_n1905_ | new_n1913_;
  assign new_n1915_ = new_n2179_ & new_n2180_ & new_n868_ & pi155 & new_n2181_;
  assign po196 = new_n1924_ | new_n1929_ | new_n1906_ | new_n1915_;
  assign new_n1917_ = new_n2179_ & new_n2180_ & new_n868_ & pi156 & new_n2181_;
  assign po197 = new_n1925_ | new_n1930_ | new_n1907_ | new_n1917_;
  assign new_n1919_ = new_n2179_ & new_n2180_ & new_n868_ & pi151 & new_n2181_;
  assign po198 = new_n1926_ | new_n1931_ | new_n1908_ | new_n1919_;
  assign new_n1921_ = new_n2182_ & new_n875_ & new_n2183_ & pi217 & new_n2184_;
  assign new_n1922_ = new_n2182_ & new_n875_ & new_n2183_ & pi218 & new_n2184_;
  assign new_n1923_ = new_n2182_ & new_n875_ & new_n2183_ & pi219 & new_n2184_;
  assign new_n1924_ = new_n2182_ & new_n875_ & new_n2183_ & pi220 & new_n2184_;
  assign new_n1925_ = new_n2182_ & new_n875_ & new_n2183_ & pi221 & new_n2184_;
  assign new_n1926_ = new_n2182_ & new_n875_ & new_n2183_ & pi222 & new_n2184_;
  assign new_n1927_ = new_n883_ & new_n2185_ & new_n2186_ & pi215 & new_n2187_;
  assign new_n1928_ = new_n883_ & new_n2185_ & new_n2186_ & pi214 & new_n2187_;
  assign new_n1929_ = new_n883_ & new_n2185_ & new_n2186_ & pi213 & new_n2187_;
  assign new_n1930_ = new_n883_ & new_n2185_ & new_n2186_ & pi212 & new_n2187_;
  assign new_n1931_ = new_n883_ & new_n2185_ & new_n2186_ & pi211 & new_n2187_;
  assign new_n1932_ = new_n2188_ & new_n2189_ & pi223 & new_n875_;
  assign new_n1933_ = new_n2188_ & new_n2189_ & pi224 & new_n875_;
  assign new_n1934_ = new_n2188_ & new_n2189_ & pi225 & new_n875_;
  assign new_n1935_ = new_n2188_ & new_n2189_ & pi226 & new_n875_;
  assign new_n1936_ = new_n2188_ & new_n2189_ & pi227 & new_n875_;
  assign new_n1937_ = new_n2188_ & new_n2189_ & pi228 & new_n875_;
  assign po199 = new_n2188_ & new_n2189_ & pi229 & new_n875_;
  assign new_n1939_ = new_n2188_ & new_n2189_ & pi230 & new_n875_;
  assign new_n1940_ = new_n2190_ & new_n876_ & pi231 & new_n2191_;
  assign po200 = new_n1932_ | new_n1940_;
  assign new_n1942_ = new_n2190_ & new_n876_ & pi232 & new_n2191_;
  assign po201 = new_n1933_ | new_n1942_;
  assign new_n1944_ = new_n2190_ & new_n876_ & pi233 & new_n2191_;
  assign po202 = new_n1934_ | new_n1944_;
  assign new_n1946_ = new_n2190_ & new_n876_ & pi234 & new_n2191_;
  assign po203 = new_n1935_ | new_n1946_;
  assign new_n1948_ = new_n2190_ & new_n876_ & pi235 & new_n2191_;
  assign po204 = new_n1936_ | new_n1948_;
  assign new_n1950_ = new_n2190_ & new_n876_ & pi236 & new_n2191_;
  assign po205 = new_n1937_ | new_n1950_;
  assign po206 = new_n1939_ | new_n1953_;
  assign new_n1953_ = new_n884_ & new_n2192_ & pi216 & new_n2193_;
  assign new_n1954_ = new_n2194_ & pi237 & new_n876_;
  assign new_n1955_ = new_n2194_ & pi238 & new_n876_;
  assign new_n1956_ = new_n540_ & pi239 & new_n2195_;
  assign po207 = new_n1954_ | new_n1956_;
  assign new_n1958_ = new_n540_ & pi240 & new_n2195_;
  assign po208 = new_n1955_ | new_n1958_;
  assign new_n1960_ = pi004 & new_n876_;
  assign new_n1961_ = pi205 & new_n2175_ & new_n1785_;
  assign new_n1962_ = pi241 | po166;
  assign new_n1963_ = ~new_n1960_;
  assign new_n1964_ = ~new_n1961_;
  assign new_n1965_ = new_n833_ & new_n1968_ & new_n1962_;
  assign new_n1966_ = pi150 & new_n1963_ & pi242 & new_n1964_;
  assign po209 = new_n1966_ | new_n1965_;
  assign new_n1968_ = ~pi242;
  assign new_n1969_ = ~pi010;
  assign new_n1970_ = ~pi011;
  assign new_n1971_ = new_n1970_ & new_n1969_;
  assign new_n1972_ = pi011 & new_n1969_;
  assign new_n1973_ = ~new_n2893_;
  assign new_n1974_ = ~new_n1972_;
  assign new_n1975_ = new_n835_ | new_n833_;
  assign new_n1976_ = pi078 & new_n828_ & new_n1975_;
  assign new_n1977_ = new_n858_ & new_n828_ & pi078;
  assign new_n1978_ = ~new_n1678_;
  assign new_n1979_ = new_n1777_ & new_n1978_ & new_n1680_ & new_n1975_ & new_n496_;
  assign new_n1980_ = new_n1777_ & new_n1978_ & new_n1680_ & new_n858_ & new_n496_;
  assign new_n1981_ = new_n1976_ | new_n1979_;
  assign new_n1982_ = new_n1980_ | new_n1977_;
  assign new_n1983_ = ~pi109;
  assign new_n1984_ = new_n2196_ & new_n2002_ & new_n1990_ & new_n2006_;
  assign new_n1985_ = new_n2196_ & new_n2002_ & new_n2903_ & new_n2006_;
  assign new_n1986_ = new_n2197_ & new_n2012_ & pi243 & new_n2013_;
  assign po210 = new_n1984_ | new_n1986_;
  assign new_n1988_ = new_n2197_ & new_n2012_ & pi244 & new_n2013_;
  assign po211 = new_n1985_ | new_n1988_;
  assign new_n1990_ = ~pi243;
  assign new_n1991_ = pi017 & pi171 & pi177;
  assign new_n1992_ = new_n936_ & new_n1771_ & new_n1510_ & pi191;
  assign new_n1993_ = new_n1509_ & new_n783_ & pi245 & new_n936_ & pi191 & new_n1771_;
  assign new_n1994_ = ~new_n1992_;
  assign new_n1995_ = new_n1766_ | new_n1991_ | new_n1764_ | pi021 | new_n1767_ | new_n1765_;
  assign new_n1996_ = new_n2007_ & new_n936_ & pi200 & new_n2000_ & new_n1510_;
  assign new_n1997_ = new_n1509_ & new_n783_ & pi245 & new_n936_ & pi200 & pi243 & pi244;
  assign new_n1998_ = new_n1992_ | new_n1997_ | new_n1996_ | new_n1993_ | new_n1995_;
  assign new_n1999_ = new_n2003_ & pi004;
  assign new_n2000_ = ~new_n1999_;
  assign new_n2001_ = new_n936_ & new_n1509_;
  assign new_n2002_ = new_n782_ & new_n1795_ & pi023;
  assign new_n2003_ = new_n860_ | new_n902_;
  assign new_n2004_ = ~new_n2001_;
  assign new_n2005_ = po065 & new_n2003_;
  assign new_n2006_ = ~new_n2005_;
  assign new_n2007_ = new_n859_ | new_n2003_;
  assign new_n2008_ = new_n2020_ & new_n2004_ & new_n2003_ & new_n1994_ & new_n2018_;
  assign new_n2009_ = new_n1761_ & new_n859_ & new_n936_ & new_n1510_ & new_n1994_ & new_n2020_;
  assign new_n2010_ = pi243 & pi244 & new_n1509_ & new_n1761_ & new_n2002_;
  assign new_n2011_ = new_n2007_ & new_n936_ & new_n1510_;
  assign new_n2012_ = ~new_n2005_;
  assign new_n2013_ = ~new_n2002_;
  assign new_n2014_ = new_n2009_ | new_n2010_ | new_n2008_;
  assign new_n2015_ = new_n2011_ | new_n2010_;
  assign new_n2016_ = ~new_n2014_;
  assign new_n2017_ = new_n936_ & new_n1755_;
  assign new_n2018_ = ~new_n2017_;
  assign new_n2019_ = new_n936_ & pi012;
  assign new_n2020_ = ~new_n2019_;
  assign new_n2021_ = new_n1851_ & new_n1974_;
  assign new_n2022_ = new_n1853_ & new_n2021_;
  assign new_n2023_ = new_n1973_ & new_n2021_;
  assign new_n2024_ = new_n1973_ & new_n1853_;
  assign new_n2025_ = new_n2023_ | new_n2024_ | new_n2022_;
  assign new_n2026_ = new_n1849_ & new_n2025_;
  assign new_n2027_ = new_n1971_ & new_n2025_;
  assign new_n2028_ = new_n1971_ & new_n1849_;
  assign new_n2029_ = new_n2027_ | new_n2028_ | new_n2026_;
  assign new_n2030_ = ~new_n2908_;
  assign new_n2031_ = ~new_n2923_;
  assign new_n2032_ = ~new_n2928_;
  assign new_n2033_ = new_n2031_ & new_n2030_;
  assign new_n2034_ = new_n2032_ & new_n2033_;
  assign new_n2035_ = ~new_n2030_;
  assign new_n2036_ = ~new_n2938_;
  assign new_n2037_ = ~new_n2943_;
  assign new_n2038_ = new_n2036_ & new_n2035_;
  assign new_n2039_ = new_n2037_ & new_n2038_;
  assign new_n2040_ = new_n2198_ & new_n2933_ & new_n1853_;
  assign new_n2041_ = new_n1867_ & new_n2963_ & new_n2199_;
  assign new_n2042_ = new_n2040_ | new_n2041_;
  assign new_n2043_ = new_n2200_ & new_n2928_ & new_n1853_;
  assign new_n2044_ = new_n1867_ & new_n2958_ & new_n2201_;
  assign new_n2045_ = new_n2043_ | new_n2044_;
  assign new_n2046_ = new_n2202_ & new_n2923_ & new_n1853_;
  assign new_n2047_ = new_n1867_ & new_n2953_ & new_n2203_;
  assign new_n2048_ = new_n2046_ | new_n2047_;
  assign new_n2049_ = new_n2204_ & new_n2908_ & new_n1853_;
  assign new_n2050_ = new_n1867_ & new_n2035_ & new_n2205_;
  assign new_n2051_ = new_n2049_ | new_n2050_;
  assign new_n2052_ = ~new_n2051_;
  assign new_n2053_ = ~new_n2048_;
  assign new_n2054_ = ~new_n2045_;
  assign new_n2055_ = new_n2053_ & new_n2052_;
  assign new_n2056_ = new_n2054_ & new_n2055_;
  assign new_n2057_ = new_n2206_ & new_n2933_ & new_n1851_;
  assign new_n2058_ = new_n1866_ & new_n2978_ & new_n2207_;
  assign new_n2059_ = new_n2057_ | new_n2058_;
  assign new_n2060_ = new_n2208_ & new_n2928_ & new_n1851_;
  assign new_n2061_ = new_n1866_ & new_n2973_ & new_n2209_;
  assign new_n2062_ = new_n2060_ | new_n2061_;
  assign new_n2063_ = new_n2210_ & new_n2923_ & new_n1851_;
  assign new_n2064_ = new_n1866_ & new_n2968_ & new_n2211_;
  assign new_n2065_ = new_n2063_ | new_n2064_;
  assign new_n2066_ = new_n2212_ & new_n2908_ & new_n1851_;
  assign new_n2067_ = new_n1866_ & new_n2052_ & new_n2213_;
  assign new_n2068_ = new_n2066_ | new_n2067_;
  assign new_n2069_ = ~new_n1871_;
  assign new_n2070_ = ~new_n1861_;
  assign new_n2071_ = ~new_n1871_;
  assign new_n2072_ = ~new_n1861_;
  assign new_n2073_ = ~new_n1871_;
  assign new_n2074_ = ~new_n1861_;
  assign new_n2075_ = ~new_n1871_;
  assign new_n2076_ = ~new_n1861_;
  assign new_n2077_ = ~new_n1870_;
  assign new_n2078_ = ~new_n1859_;
  assign new_n2079_ = ~new_n1870_;
  assign new_n2080_ = ~new_n1859_;
  assign new_n2081_ = ~new_n1870_;
  assign new_n2082_ = ~new_n1859_;
  assign new_n2083_ = ~new_n1870_;
  assign new_n2084_ = ~new_n1859_;
  assign new_n2085_ = ~new_n902_ | ~po065;
  assign new_n2086_ = ~new_n2015_;
  assign new_n2087_ = ~new_n902_ | ~po065;
  assign new_n2088_ = ~new_n860_ | ~po065;
  assign new_n2089_ = ~new_n2015_;
  assign new_n2090_ = ~new_n860_ | ~po065;
  assign new_n2091_ = ~new_n2007_;
  assign new_n2092_ = ~new_n1459_;
  assign new_n2093_ = ~new_n2007_;
  assign new_n2094_ = ~new_n1459_;
  assign new_n2095_ = ~new_n1485_;
  assign new_n2096_ = ~new_n1072_ | ~new_n860_ | ~new_n1510_;
  assign new_n2097_ = ~new_n1072_ | ~new_n860_ | ~new_n1510_;
  assign new_n2098_ = ~new_n1715_;
  assign new_n2099_ = ~new_n1485_;
  assign new_n2100_ = ~new_n1072_ | ~new_n860_ | ~new_n1510_;
  assign new_n2101_ = ~new_n1485_;
  assign new_n2102_ = ~new_n1715_;
  assign new_n2103_ = ~new_n1072_ | ~new_n860_ | ~new_n1510_;
  assign new_n2104_ = ~new_n1715_;
  assign new_n2105_ = ~new_n1472_;
  assign new_n2106_ = new_n2105_ & new_n1466_;
  assign new_n2107_ = ~new_n1466_;
  assign new_n2108_ = ~new_n1209_;
  assign new_n2109_ = ~new_n1210_;
  assign new_n2110_ = ~new_n1209_;
  assign new_n2111_ = ~new_n1210_;
  assign new_n2112_ = ~new_n1481_;
  assign new_n2113_ = ~new_n1486_;
  assign new_n2114_ = ~new_n1481_;
  assign new_n2115_ = ~new_n1486_;
  assign new_n2116_ = ~new_n1481_;
  assign new_n2117_ = ~new_n1486_;
  assign new_n2118_ = ~new_n1982_;
  assign new_n2119_ = ~new_n1362_;
  assign new_n2120_ = ~new_n1977_;
  assign new_n2121_ = ~new_n1366_;
  assign new_n2122_ = ~new_n1869_;
  assign new_n2123_ = ~new_n1857_;
  assign new_n2124_ = ~new_n1869_;
  assign new_n2125_ = ~new_n1857_;
  assign new_n2126_ = ~new_n1869_;
  assign new_n2127_ = ~new_n1857_;
  assign new_n2128_ = ~new_n1869_;
  assign new_n2129_ = ~new_n1857_;
  assign new_n2130_ = ~new_n1868_;
  assign new_n2131_ = ~new_n1855_;
  assign new_n2132_ = ~new_n1868_;
  assign new_n2133_ = ~new_n1855_;
  assign new_n2134_ = ~new_n1868_;
  assign new_n2135_ = ~new_n1855_;
  assign new_n2136_ = ~new_n1868_;
  assign new_n2137_ = ~new_n1855_;
  assign new_n2138_ = ~new_n537_;
  assign new_n2139_ = ~new_n854_ | ~new_n936_;
  assign new_n2140_ = ~new_n1981_;
  assign new_n2141_ = ~new_n1724_;
  assign new_n2142_ = ~new_n1976_;
  assign new_n2143_ = ~new_n1728_;
  assign new_n2144_ = ~new_n1795_;
  assign new_n2145_ = ~pi065;
  assign new_n2146_ = ~pi066;
  assign new_n2147_ = ~new_n878_;
  assign new_n2148_ = ~pi244;
  assign new_n2149_ = ~pi243;
  assign new_n2150_ = ~new_n878_;
  assign new_n2151_ = ~po071;
  assign new_n2152_ = ~po070;
  assign new_n2153_ = ~new_n1795_;
  assign new_n2154_ = ~pi246;
  assign new_n2155_ = ~pi247;
  assign new_n2156_ = ~new_n594_;
  assign new_n2157_ = ~po090;
  assign new_n2158_ = ~po089;
  assign new_n2159_ = ~po088;
  assign new_n2160_ = ~po087;
  assign new_n2161_ = ~po086;
  assign new_n2162_ = ~po085;
  assign new_n2163_ = ~po084;
  assign new_n2164_ = ~po083;
  assign new_n2165_ = ~po082;
  assign new_n2166_ = ~pi022;
  assign new_n2167_ = ~po077;
  assign new_n2168_ = ~po076;
  assign new_n2169_ = ~po075;
  assign new_n2170_ = ~po074;
  assign new_n2171_ = ~po073;
  assign new_n2172_ = ~po072;
  assign new_n2173_ = ~po071;
  assign new_n2174_ = ~po070;
  assign new_n2175_ = ~pi215;
  assign new_n2176_ = ~new_n883_;
  assign new_n2177_ = ~new_n875_;
  assign new_n2178_ = ~new_n868_;
  assign new_n2179_ = ~new_n883_;
  assign new_n2180_ = ~new_n875_;
  assign new_n2181_ = ~new_n869_;
  assign new_n2182_ = ~new_n883_;
  assign new_n2183_ = ~new_n868_;
  assign new_n2184_ = ~new_n869_;
  assign new_n2185_ = ~new_n875_;
  assign new_n2186_ = ~new_n868_;
  assign new_n2187_ = ~new_n869_;
  assign new_n2188_ = ~new_n884_;
  assign new_n2189_ = ~new_n876_;
  assign new_n2190_ = ~new_n884_;
  assign new_n2191_ = ~new_n875_;
  assign new_n2192_ = ~new_n876_;
  assign new_n2193_ = ~new_n875_;
  assign new_n2194_ = ~new_n540_;
  assign new_n2195_ = ~new_n876_;
  assign new_n2196_ = ~new_n2012_ | ~new_n2013_;
  assign new_n2197_ = ~new_n2002_ | ~new_n2006_;
  assign new_n2198_ = ~new_n1867_;
  assign new_n2199_ = ~new_n1853_;
  assign new_n2200_ = ~new_n1867_;
  assign new_n2201_ = ~new_n1853_;
  assign new_n2202_ = ~new_n1867_;
  assign new_n2203_ = ~new_n1853_;
  assign new_n2204_ = ~new_n1867_;
  assign new_n2205_ = ~new_n1853_;
  assign new_n2206_ = ~new_n1866_;
  assign new_n2207_ = ~new_n1851_;
  assign new_n2208_ = ~new_n1866_;
  assign new_n2209_ = ~new_n1851_;
  assign new_n2210_ = ~new_n1866_;
  assign new_n2211_ = ~new_n1851_;
  assign new_n2212_ = ~new_n1866_;
  assign new_n2213_ = ~new_n1851_;
  assign new_n2214_ = ~new_n2258_;
  assign new_n2215_ = ~pi000;
  assign new_n2216_ = new_n2258_ & new_n2215_;
  assign new_n2217_ = new_n2214_ & pi000;
  assign new_n2218_ = new_n2216_ | new_n2217_;
  assign new_n2219_ = ~new_n2253_;
  assign new_n2220_ = ~pi001;
  assign new_n2221_ = new_n2253_ & new_n2220_;
  assign new_n2222_ = new_n2219_ & pi001;
  assign new_n2223_ = new_n2221_ | new_n2222_;
  assign new_n2224_ = ~new_n2248_;
  assign new_n2225_ = ~pi002;
  assign new_n2226_ = new_n2248_ & new_n2225_;
  assign new_n2227_ = new_n2224_ & pi002;
  assign new_n2228_ = new_n2226_ | new_n2227_;
  assign new_n2229_ = ~new_n1859_;
  assign new_n2230_ = ~new_n2598_;
  assign new_n2231_ = new_n1859_ & new_n2230_;
  assign new_n2232_ = new_n2229_ & new_n2598_;
  assign new_n2233_ = new_n2231_ | new_n2232_;
  assign new_n2234_ = ~new_n1861_;
  assign new_n2235_ = ~new_n2613_;
  assign new_n2236_ = new_n1861_ & new_n2235_;
  assign new_n2237_ = new_n2234_ & new_n2613_;
  assign new_n2238_ = new_n2236_ | new_n2237_;
  assign new_n2239_ = ~new_n1847_;
  assign new_n2240_ = ~new_n2618_;
  assign new_n2241_ = new_n1847_ & new_n2240_;
  assign new_n2242_ = new_n2239_ & new_n2618_;
  assign new_n2243_ = new_n2241_ | new_n2242_;
  assign new_n2244_ = ~new_n2238_;
  assign new_n2245_ = ~new_n595_;
  assign new_n2246_ = new_n2238_ & new_n2245_;
  assign new_n2247_ = new_n2244_ & new_n595_;
  assign new_n2248_ = new_n2246_ | new_n2247_;
  assign new_n2249_ = ~new_n599_;
  assign new_n2250_ = ~new_n2243_;
  assign new_n2251_ = new_n599_ & new_n2250_;
  assign new_n2252_ = new_n2249_ & new_n2243_;
  assign new_n2253_ = new_n2251_ | new_n2252_;
  assign new_n2254_ = ~new_n2623_;
  assign new_n2255_ = ~new_n603_;
  assign new_n2256_ = new_n2623_ & new_n2255_;
  assign new_n2257_ = new_n2254_ & new_n603_;
  assign new_n2258_ = new_n2256_ | new_n2257_;
  assign new_n2259_ = ~new_n2248_;
  assign new_n2260_ = ~new_n491_;
  assign new_n2261_ = new_n2248_ & new_n2260_;
  assign new_n2262_ = new_n2259_ & new_n491_;
  assign new_n2263_ = new_n2261_ | new_n2262_;
  assign new_n2264_ = ~new_n2253_;
  assign new_n2265_ = ~new_n604_;
  assign new_n2266_ = new_n2253_ & new_n2265_;
  assign new_n2267_ = new_n2264_ & new_n604_;
  assign new_n2268_ = new_n2266_ | new_n2267_;
  assign new_n2269_ = ~new_n2258_;
  assign new_n2270_ = ~new_n605_;
  assign new_n2271_ = new_n2258_ & new_n2270_;
  assign new_n2272_ = new_n2269_ & new_n605_;
  assign new_n2273_ = new_n2271_ | new_n2272_;
  assign new_n2274_ = ~new_n2263_;
  assign new_n2275_ = ~new_n606_;
  assign new_n2276_ = new_n2263_ & new_n2275_;
  assign new_n2277_ = new_n2274_ & new_n606_;
  assign new_n2278_ = new_n2276_ | new_n2277_;
  assign new_n2279_ = ~new_n2268_;
  assign new_n2280_ = ~new_n609_;
  assign new_n2281_ = new_n2268_ & new_n2280_;
  assign new_n2282_ = new_n2279_ & new_n609_;
  assign new_n2283_ = new_n2281_ | new_n2282_;
  assign new_n2284_ = ~new_n2273_;
  assign new_n2285_ = ~new_n610_;
  assign new_n2286_ = new_n2273_ & new_n2285_;
  assign new_n2287_ = new_n2284_ & new_n610_;
  assign new_n2288_ = new_n2286_ | new_n2287_;
  assign new_n2289_ = ~new_n619_;
  assign new_n2290_ = ~new_n623_;
  assign new_n2291_ = new_n619_ & new_n2290_;
  assign new_n2292_ = new_n2289_ & new_n623_;
  assign new_n2293_ = new_n2291_ | new_n2292_;
  assign new_n2294_ = ~new_n616_;
  assign new_n2295_ = ~new_n626_;
  assign new_n2296_ = new_n616_ & new_n2295_;
  assign new_n2297_ = new_n2294_ & new_n626_;
  assign new_n2298_ = new_n2296_ | new_n2297_;
  assign new_n2299_ = ~new_n613_;
  assign new_n2300_ = ~new_n627_;
  assign new_n2301_ = new_n613_ & new_n2300_;
  assign new_n2302_ = new_n2299_ & new_n627_;
  assign new_n2303_ = new_n2301_ | new_n2302_;
  assign new_n2304_ = ~pi248;
  assign new_n2305_ = ~pi249;
  assign new_n2306_ = pi248 & new_n2305_;
  assign new_n2307_ = new_n2304_ & pi249;
  assign new_n2308_ = new_n2306_ | new_n2307_;
  assign new_n2309_ = ~pi250;
  assign new_n2310_ = ~pi251;
  assign new_n2311_ = pi250 & new_n2310_;
  assign new_n2312_ = new_n2309_ & pi251;
  assign new_n2313_ = new_n2311_ | new_n2312_;
  assign new_n2314_ = ~pi252;
  assign new_n2315_ = ~pi025;
  assign new_n2316_ = pi252 & new_n2315_;
  assign new_n2317_ = new_n2314_ & pi025;
  assign new_n2318_ = new_n2316_ | new_n2317_;
  assign new_n2319_ = ~pi129;
  assign new_n2320_ = ~new_n784_;
  assign new_n2321_ = pi129 & new_n2320_;
  assign new_n2322_ = new_n2319_ & new_n784_;
  assign po212 = new_n2321_ | new_n2322_;
  assign new_n2324_ = ~pi048;
  assign new_n2325_ = ~new_n785_;
  assign new_n2326_ = pi048 & new_n2325_;
  assign new_n2327_ = new_n2324_ & new_n785_;
  assign po213 = new_n2326_ | new_n2327_;
  assign new_n2329_ = ~pi049;
  assign new_n2330_ = ~new_n786_;
  assign new_n2331_ = pi049 & new_n2330_;
  assign new_n2332_ = new_n2329_ & new_n786_;
  assign po214 = new_n2331_ | new_n2332_;
  assign new_n2334_ = ~pi047;
  assign new_n2335_ = ~new_n787_;
  assign new_n2336_ = pi047 & new_n2335_;
  assign new_n2337_ = new_n2334_ & new_n787_;
  assign po215 = new_n2336_ | new_n2337_;
  assign new_n2339_ = ~pi050;
  assign new_n2340_ = ~new_n788_;
  assign new_n2341_ = pi050 & new_n2340_;
  assign new_n2342_ = new_n2339_ & new_n788_;
  assign po216 = new_n2341_ | new_n2342_;
  assign new_n2344_ = ~pi046;
  assign new_n2345_ = ~new_n789_;
  assign new_n2346_ = pi046 & new_n2345_;
  assign new_n2347_ = new_n2344_ & new_n789_;
  assign po217 = new_n2346_ | new_n2347_;
  assign new_n2349_ = ~pi051;
  assign new_n2350_ = ~pi045;
  assign new_n2351_ = pi051 & new_n2350_;
  assign new_n2352_ = new_n2349_ & pi045;
  assign po218 = new_n2351_ | new_n2352_;
  assign new_n2354_ = ~new_n2059_;
  assign new_n2355_ = ~new_n1339_;
  assign new_n2356_ = new_n2059_ & new_n2355_;
  assign new_n2357_ = new_n2354_ & new_n1339_;
  assign new_n2358_ = new_n2356_ | new_n2357_;
  assign new_n2359_ = ~new_n2062_;
  assign new_n2360_ = ~new_n1337_;
  assign new_n2361_ = new_n2062_ & new_n2360_;
  assign new_n2362_ = new_n2359_ & new_n1337_;
  assign new_n2363_ = new_n2361_ | new_n2362_;
  assign new_n2364_ = ~new_n2065_;
  assign new_n2365_ = ~new_n1335_;
  assign new_n2366_ = new_n2065_ & new_n2365_;
  assign new_n2367_ = new_n2364_ & new_n1335_;
  assign new_n2368_ = new_n2366_ | new_n2367_;
  assign new_n2369_ = ~new_n2068_;
  assign new_n2370_ = ~new_n1333_;
  assign new_n2371_ = new_n2068_ & new_n2370_;
  assign new_n2372_ = new_n2369_ & new_n1333_;
  assign new_n2373_ = new_n2371_ | new_n2372_;
  assign new_n2374_ = ~new_n2042_;
  assign new_n2375_ = ~new_n1339_;
  assign new_n2376_ = new_n2042_ & new_n2375_;
  assign new_n2377_ = new_n2374_ & new_n1339_;
  assign new_n2378_ = new_n2376_ | new_n2377_;
  assign new_n2379_ = ~new_n2045_;
  assign new_n2380_ = ~new_n1337_;
  assign new_n2381_ = new_n2045_ & new_n2380_;
  assign new_n2382_ = new_n2379_ & new_n1337_;
  assign new_n2383_ = new_n2381_ | new_n2382_;
  assign new_n2384_ = ~new_n2048_;
  assign new_n2385_ = ~new_n1335_;
  assign new_n2386_ = new_n2048_ & new_n2385_;
  assign new_n2387_ = new_n2384_ & new_n1335_;
  assign new_n2388_ = new_n2386_ | new_n2387_;
  assign new_n2389_ = ~new_n2051_;
  assign new_n2390_ = ~new_n1333_;
  assign new_n2391_ = new_n2051_ & new_n2390_;
  assign new_n2392_ = new_n2389_ & new_n1333_;
  assign new_n2393_ = new_n2391_ | new_n2392_;
  assign new_n2394_ = ~new_n2948_;
  assign new_n2395_ = ~new_n1339_;
  assign new_n2396_ = new_n2948_ & new_n2395_;
  assign new_n2397_ = new_n2394_ & new_n1339_;
  assign new_n2398_ = new_n2396_ | new_n2397_;
  assign new_n2399_ = ~new_n2943_;
  assign new_n2400_ = ~new_n1337_;
  assign new_n2401_ = new_n2943_ & new_n2400_;
  assign new_n2402_ = new_n2399_ & new_n1337_;
  assign new_n2403_ = new_n2401_ | new_n2402_;
  assign new_n2404_ = ~new_n2938_;
  assign new_n2405_ = ~new_n1335_;
  assign new_n2406_ = new_n2938_ & new_n2405_;
  assign new_n2407_ = new_n2404_ & new_n1335_;
  assign new_n2408_ = new_n2406_ | new_n2407_;
  assign new_n2409_ = ~new_n2030_;
  assign new_n2410_ = ~new_n1333_;
  assign new_n2411_ = new_n2030_ & new_n2410_;
  assign new_n2412_ = new_n2409_ & new_n1333_;
  assign new_n2413_ = new_n2411_ | new_n2412_;
  assign new_n2414_ = ~new_n2933_;
  assign new_n2415_ = ~new_n1339_;
  assign new_n2416_ = new_n2933_ & new_n2415_;
  assign new_n2417_ = new_n2414_ & new_n1339_;
  assign new_n2418_ = new_n2416_ | new_n2417_;
  assign new_n2419_ = ~new_n2928_;
  assign new_n2420_ = ~new_n1337_;
  assign new_n2421_ = new_n2928_ & new_n2420_;
  assign new_n2422_ = new_n2419_ & new_n1337_;
  assign new_n2423_ = new_n2421_ | new_n2422_;
  assign new_n2424_ = ~new_n2923_;
  assign new_n2425_ = ~new_n1335_;
  assign new_n2426_ = new_n2923_ & new_n2425_;
  assign new_n2427_ = new_n2424_ & new_n1335_;
  assign new_n2428_ = new_n2426_ | new_n2427_;
  assign new_n2429_ = ~new_n2908_;
  assign new_n2430_ = ~new_n1333_;
  assign new_n2431_ = new_n2908_ & new_n2430_;
  assign new_n2432_ = new_n2429_ & new_n1333_;
  assign new_n2433_ = new_n2431_ | new_n2432_;
  assign new_n2434_ = ~new_n1420_;
  assign new_n2435_ = ~new_n1339_;
  assign new_n2436_ = new_n1420_ & new_n2435_;
  assign new_n2437_ = new_n2434_ & new_n1339_;
  assign new_n2438_ = new_n2436_ | new_n2437_;
  assign new_n2439_ = ~new_n1423_;
  assign new_n2440_ = ~new_n1337_;
  assign new_n2441_ = new_n1423_ & new_n2440_;
  assign new_n2442_ = new_n2439_ & new_n1337_;
  assign new_n2443_ = new_n2441_ | new_n2442_;
  assign new_n2444_ = ~new_n1426_;
  assign new_n2445_ = ~new_n1335_;
  assign new_n2446_ = new_n1426_ & new_n2445_;
  assign new_n2447_ = new_n2444_ & new_n1335_;
  assign new_n2448_ = new_n2446_ | new_n2447_;
  assign new_n2449_ = ~new_n1429_;
  assign new_n2450_ = ~new_n1333_;
  assign new_n2451_ = new_n1429_ & new_n2450_;
  assign new_n2452_ = new_n2449_ & new_n1333_;
  assign new_n2453_ = new_n2451_ | new_n2452_;
  assign new_n2454_ = ~new_n1403_;
  assign new_n2455_ = ~new_n1339_;
  assign new_n2456_ = new_n1403_ & new_n2455_;
  assign new_n2457_ = new_n2454_ & new_n1339_;
  assign new_n2458_ = new_n2456_ | new_n2457_;
  assign new_n2459_ = ~new_n1406_;
  assign new_n2460_ = ~new_n1337_;
  assign new_n2461_ = new_n1406_ & new_n2460_;
  assign new_n2462_ = new_n2459_ & new_n1337_;
  assign new_n2463_ = new_n2461_ | new_n2462_;
  assign new_n2464_ = ~new_n1409_;
  assign new_n2465_ = ~new_n1335_;
  assign new_n2466_ = new_n1409_ & new_n2465_;
  assign new_n2467_ = new_n2464_ & new_n1335_;
  assign new_n2468_ = new_n2466_ | new_n2467_;
  assign new_n2469_ = ~new_n1412_;
  assign new_n2470_ = ~new_n1333_;
  assign new_n2471_ = new_n1412_ & new_n2470_;
  assign new_n2472_ = new_n2469_ & new_n1333_;
  assign new_n2473_ = new_n2471_ | new_n2472_;
  assign new_n2474_ = ~new_n2638_;
  assign new_n2475_ = ~new_n1339_;
  assign new_n2476_ = new_n2638_ & new_n2475_;
  assign new_n2477_ = new_n2474_ & new_n1339_;
  assign new_n2478_ = new_n2476_ | new_n2477_;
  assign new_n2479_ = ~new_n2633_;
  assign new_n2480_ = ~new_n1337_;
  assign new_n2481_ = new_n2633_ & new_n2480_;
  assign new_n2482_ = new_n2479_ & new_n1337_;
  assign new_n2483_ = new_n2481_ | new_n2482_;
  assign new_n2484_ = ~new_n2628_;
  assign new_n2485_ = ~new_n1335_;
  assign new_n2486_ = new_n2628_ & new_n2485_;
  assign new_n2487_ = new_n2484_ & new_n1335_;
  assign new_n2488_ = new_n2486_ | new_n2487_;
  assign new_n2489_ = ~new_n1391_;
  assign new_n2490_ = ~new_n1333_;
  assign new_n2491_ = new_n1391_ & new_n2490_;
  assign new_n2492_ = new_n2489_ & new_n1333_;
  assign new_n2493_ = new_n2491_ | new_n2492_;
  assign new_n2494_ = ~new_n2623_;
  assign new_n2495_ = ~new_n1339_;
  assign new_n2496_ = new_n2623_ & new_n2495_;
  assign new_n2497_ = new_n2494_ & new_n1339_;
  assign new_n2498_ = new_n2496_ | new_n2497_;
  assign new_n2499_ = ~new_n2618_;
  assign new_n2500_ = ~new_n1337_;
  assign new_n2501_ = new_n2618_ & new_n2500_;
  assign new_n2502_ = new_n2499_ & new_n1337_;
  assign new_n2503_ = new_n2501_ | new_n2502_;
  assign new_n2504_ = ~new_n2613_;
  assign new_n2505_ = ~new_n1335_;
  assign new_n2506_ = new_n2613_ & new_n2505_;
  assign new_n2507_ = new_n2504_ & new_n1335_;
  assign new_n2508_ = new_n2506_ | new_n2507_;
  assign new_n2509_ = ~new_n2598_;
  assign new_n2510_ = ~new_n1333_;
  assign new_n2511_ = new_n2598_ & new_n2510_;
  assign new_n2512_ = new_n2509_ & new_n1333_;
  assign new_n2513_ = new_n2511_ | new_n2512_;
  assign new_n2514_ = ~new_n630_;
  assign new_n2515_ = ~new_n1339_;
  assign new_n2516_ = new_n630_ & new_n2515_;
  assign new_n2517_ = new_n2514_ & new_n1339_;
  assign new_n2518_ = new_n2516_ | new_n2517_;
  assign new_n2519_ = ~new_n633_;
  assign new_n2520_ = ~new_n1337_;
  assign new_n2521_ = new_n633_ & new_n2520_;
  assign new_n2522_ = new_n2519_ & new_n1337_;
  assign new_n2523_ = new_n2521_ | new_n2522_;
  assign new_n2524_ = ~new_n636_;
  assign new_n2525_ = ~new_n1335_;
  assign new_n2526_ = new_n636_ & new_n2525_;
  assign new_n2527_ = new_n2524_ & new_n1335_;
  assign new_n2528_ = new_n2526_ | new_n2527_;
  assign new_n2529_ = ~new_n639_;
  assign new_n2530_ = ~new_n1333_;
  assign new_n2531_ = new_n639_ & new_n2530_;
  assign new_n2532_ = new_n2529_ & new_n1333_;
  assign new_n2533_ = new_n2531_ | new_n2532_;
  assign new_n2534_ = ~new_n613_;
  assign new_n2535_ = ~new_n1339_;
  assign new_n2536_ = new_n613_ & new_n2535_;
  assign new_n2537_ = new_n2534_ & new_n1339_;
  assign new_n2538_ = new_n2536_ | new_n2537_;
  assign new_n2539_ = ~new_n616_;
  assign new_n2540_ = ~new_n1337_;
  assign new_n2541_ = new_n616_ & new_n2540_;
  assign new_n2542_ = new_n2539_ & new_n1337_;
  assign new_n2543_ = new_n2541_ | new_n2542_;
  assign new_n2544_ = ~new_n619_;
  assign new_n2545_ = ~new_n1335_;
  assign new_n2546_ = new_n619_ & new_n2545_;
  assign new_n2547_ = new_n2544_ & new_n1335_;
  assign new_n2548_ = new_n2546_ | new_n2547_;
  assign new_n2549_ = ~new_n622_;
  assign new_n2550_ = ~new_n1333_;
  assign new_n2551_ = new_n622_ & new_n2550_;
  assign new_n2552_ = new_n2549_ & new_n1333_;
  assign new_n2553_ = new_n2551_ | new_n2552_;
  assign new_n2554_ = ~new_n2273_;
  assign new_n2555_ = ~new_n1339_;
  assign new_n2556_ = new_n2273_ & new_n2555_;
  assign new_n2557_ = new_n2554_ & new_n1339_;
  assign new_n2558_ = new_n2556_ | new_n2557_;
  assign new_n2559_ = ~new_n2268_;
  assign new_n2560_ = ~new_n1337_;
  assign new_n2561_ = new_n2268_ & new_n2560_;
  assign new_n2562_ = new_n2559_ & new_n1337_;
  assign new_n2563_ = new_n2561_ | new_n2562_;
  assign new_n2564_ = ~new_n2263_;
  assign new_n2565_ = ~new_n1335_;
  assign new_n2566_ = new_n2263_ & new_n2565_;
  assign new_n2567_ = new_n2564_ & new_n1335_;
  assign new_n2568_ = new_n2566_ | new_n2567_;
  assign new_n2569_ = ~new_n491_;
  assign new_n2570_ = ~new_n1333_;
  assign new_n2571_ = new_n491_ & new_n2570_;
  assign new_n2572_ = new_n2569_ & new_n1333_;
  assign new_n2573_ = new_n2571_ | new_n2572_;
  assign new_n2574_ = ~new_n2258_;
  assign new_n2575_ = ~new_n1339_;
  assign new_n2576_ = new_n2258_ & new_n2575_;
  assign new_n2577_ = new_n2574_ & new_n1339_;
  assign new_n2578_ = new_n2576_ | new_n2577_;
  assign new_n2579_ = ~new_n2253_;
  assign new_n2580_ = ~new_n1337_;
  assign new_n2581_ = new_n2253_ & new_n2580_;
  assign new_n2582_ = new_n2579_ & new_n1337_;
  assign new_n2583_ = new_n2581_ | new_n2582_;
  assign new_n2584_ = ~new_n2248_;
  assign new_n2585_ = ~new_n1335_;
  assign new_n2586_ = new_n2248_ & new_n2585_;
  assign new_n2587_ = new_n2584_ & new_n1335_;
  assign new_n2588_ = new_n2586_ | new_n2587_;
  assign new_n2589_ = ~new_n2233_;
  assign new_n2590_ = ~new_n1333_;
  assign new_n2591_ = new_n2233_ & new_n2590_;
  assign new_n2592_ = new_n2589_ & new_n1333_;
  assign new_n2593_ = new_n2591_ | new_n2592_;
  assign new_n2594_ = ~new_n1855_;
  assign new_n2595_ = ~new_n2908_;
  assign new_n2596_ = new_n1855_ & new_n2595_;
  assign new_n2597_ = new_n2594_ & new_n2908_;
  assign new_n2598_ = new_n2596_ | new_n2597_;
  assign new_n2599_ = ~new_n1857_;
  assign new_n2600_ = ~new_n2923_;
  assign new_n2601_ = new_n1857_ & new_n2600_;
  assign new_n2602_ = new_n2599_ & new_n2923_;
  assign new_n2603_ = new_n2601_ | new_n2602_;
  assign new_n2604_ = ~new_n1848_;
  assign new_n2605_ = ~new_n2928_;
  assign new_n2606_ = new_n1848_ & new_n2605_;
  assign new_n2607_ = new_n2604_ & new_n2928_;
  assign new_n2608_ = new_n2606_ | new_n2607_;
  assign new_n2609_ = ~new_n2603_;
  assign new_n2610_ = ~new_n1382_;
  assign new_n2611_ = new_n2603_ & new_n2610_;
  assign new_n2612_ = new_n2609_ & new_n1382_;
  assign new_n2613_ = new_n2611_ | new_n2612_;
  assign new_n2614_ = ~new_n1386_;
  assign new_n2615_ = ~new_n2608_;
  assign new_n2616_ = new_n1386_ & new_n2615_;
  assign new_n2617_ = new_n2614_ & new_n2608_;
  assign new_n2618_ = new_n2616_ | new_n2617_;
  assign new_n2619_ = ~new_n2933_;
  assign new_n2620_ = ~new_n1390_;
  assign new_n2621_ = new_n2933_ & new_n2620_;
  assign new_n2622_ = new_n2619_ & new_n1390_;
  assign new_n2623_ = new_n2621_ | new_n2622_;
  assign new_n2624_ = ~new_n2613_;
  assign new_n2625_ = ~new_n1391_;
  assign new_n2626_ = new_n2613_ & new_n2625_;
  assign new_n2627_ = new_n2624_ & new_n1391_;
  assign new_n2628_ = new_n2626_ | new_n2627_;
  assign new_n2629_ = ~new_n2618_;
  assign new_n2630_ = ~new_n1394_;
  assign new_n2631_ = new_n2618_ & new_n2630_;
  assign new_n2632_ = new_n2629_ & new_n1394_;
  assign new_n2633_ = new_n2631_ | new_n2632_;
  assign new_n2634_ = ~new_n2623_;
  assign new_n2635_ = ~new_n1395_;
  assign new_n2636_ = new_n2623_ & new_n2635_;
  assign new_n2637_ = new_n2634_ & new_n1395_;
  assign new_n2638_ = new_n2636_ | new_n2637_;
  assign new_n2639_ = ~new_n2628_;
  assign new_n2640_ = ~new_n1396_;
  assign new_n2641_ = new_n2628_ & new_n2640_;
  assign new_n2642_ = new_n2639_ & new_n1396_;
  assign new_n2643_ = new_n2641_ | new_n2642_;
  assign new_n2644_ = ~new_n2633_;
  assign new_n2645_ = ~new_n1399_;
  assign new_n2646_ = new_n2633_ & new_n2645_;
  assign new_n2647_ = new_n2644_ & new_n1399_;
  assign new_n2648_ = new_n2646_ | new_n2647_;
  assign new_n2649_ = ~new_n2638_;
  assign new_n2650_ = ~new_n1400_;
  assign new_n2651_ = new_n2638_ & new_n2650_;
  assign new_n2652_ = new_n2649_ & new_n1400_;
  assign new_n2653_ = new_n2651_ | new_n2652_;
  assign new_n2654_ = ~new_n1409_;
  assign new_n2655_ = ~new_n1413_;
  assign new_n2656_ = new_n1409_ & new_n2655_;
  assign new_n2657_ = new_n2654_ & new_n1413_;
  assign new_n2658_ = new_n2656_ | new_n2657_;
  assign new_n2659_ = ~new_n1406_;
  assign new_n2660_ = ~new_n1416_;
  assign new_n2661_ = new_n1406_ & new_n2660_;
  assign new_n2662_ = new_n2659_ & new_n1416_;
  assign new_n2663_ = new_n2661_ | new_n2662_;
  assign new_n2664_ = ~new_n1403_;
  assign new_n2665_ = ~new_n1417_;
  assign new_n2666_ = new_n1403_ & new_n2665_;
  assign new_n2667_ = new_n2664_ & new_n1417_;
  assign new_n2668_ = new_n2666_ | new_n2667_;
  assign new_n2669_ = ~pi206;
  assign new_n2670_ = ~new_n1435_;
  assign new_n2671_ = pi206 & new_n2670_;
  assign new_n2672_ = new_n2669_ & new_n1435_;
  assign po219 = new_n2671_ | new_n2672_;
  assign new_n2674_ = ~pi159;
  assign new_n2675_ = ~new_n1436_;
  assign new_n2676_ = pi159 & new_n2675_;
  assign new_n2677_ = new_n2674_ & new_n1436_;
  assign po220 = new_n2676_ | new_n2677_;
  assign new_n2679_ = ~pi160;
  assign new_n2680_ = ~new_n1437_;
  assign new_n2681_ = pi160 & new_n2680_;
  assign new_n2682_ = new_n2679_ & new_n1437_;
  assign po221 = new_n2681_ | new_n2682_;
  assign new_n2684_ = ~pi158;
  assign new_n2685_ = ~new_n1438_;
  assign new_n2686_ = pi158 & new_n2685_;
  assign new_n2687_ = new_n2684_ & new_n1438_;
  assign po222 = new_n2686_ | new_n2687_;
  assign new_n2689_ = ~pi161;
  assign new_n2690_ = ~pi157;
  assign new_n2691_ = pi161 & new_n2690_;
  assign new_n2692_ = new_n2689_ & pi157;
  assign po223 = new_n2691_ | new_n2692_;
  assign new_n2694_ = ~pi253;
  assign new_n2695_ = ~pi254;
  assign new_n2696_ = pi253 & new_n2695_;
  assign new_n2697_ = new_n2694_ & pi254;
  assign new_n2698_ = new_n2696_ | new_n2697_;
  assign new_n2699_ = ~pi247;
  assign new_n2700_ = ~pi246;
  assign new_n2701_ = pi247 & new_n2700_;
  assign new_n2702_ = new_n2699_ & pi246;
  assign new_n2703_ = new_n2701_ | new_n2702_;
  assign new_n2704_ = ~pi146;
  assign new_n2705_ = ~pi147;
  assign new_n2706_ = pi146 & new_n2705_;
  assign new_n2707_ = new_n2704_ & pi147;
  assign new_n2708_ = new_n2706_ | new_n2707_;
  assign new_n2709_ = ~pi144;
  assign new_n2710_ = ~pi145;
  assign new_n2711_ = pi144 & new_n2710_;
  assign new_n2712_ = new_n2709_ & pi145;
  assign new_n2713_ = new_n2711_ | new_n2712_;
  assign new_n2714_ = ~pi142;
  assign new_n2715_ = ~pi143;
  assign new_n2716_ = pi142 & new_n2715_;
  assign new_n2717_ = new_n2714_ & pi143;
  assign new_n2718_ = new_n2716_ | new_n2717_;
  assign new_n2719_ = ~pi140;
  assign new_n2720_ = ~pi141;
  assign new_n2721_ = pi140 & new_n2720_;
  assign new_n2722_ = new_n2719_ & pi141;
  assign new_n2723_ = new_n2721_ | new_n2722_;
  assign new_n2724_ = ~pi138;
  assign new_n2725_ = ~pi139;
  assign new_n2726_ = pi138 & new_n2725_;
  assign new_n2727_ = new_n2724_ & pi139;
  assign new_n2728_ = new_n2726_ | new_n2727_;
  assign new_n2729_ = ~pi066;
  assign new_n2730_ = ~pi065;
  assign new_n2731_ = pi066 & new_n2730_;
  assign new_n2732_ = new_n2729_ & pi065;
  assign new_n2733_ = new_n2731_ | new_n2732_;
  assign new_n2734_ = ~new_n2703_;
  assign new_n2735_ = ~new_n2698_;
  assign new_n2736_ = new_n2703_ & new_n2735_;
  assign new_n2737_ = new_n2734_ & new_n2698_;
  assign new_n2738_ = new_n2736_ | new_n2737_;
  assign new_n2739_ = ~new_n2713_;
  assign new_n2740_ = ~new_n2708_;
  assign new_n2741_ = new_n2713_ & new_n2740_;
  assign new_n2742_ = new_n2739_ & new_n2708_;
  assign new_n2743_ = new_n2741_ | new_n2742_;
  assign new_n2744_ = ~new_n2723_;
  assign new_n2745_ = ~new_n2718_;
  assign new_n2746_ = new_n2723_ & new_n2745_;
  assign new_n2747_ = new_n2744_ & new_n2718_;
  assign new_n2748_ = new_n2746_ | new_n2747_;
  assign new_n2749_ = ~new_n2733_;
  assign new_n2750_ = ~new_n2728_;
  assign new_n2751_ = new_n2733_ & new_n2750_;
  assign new_n2752_ = new_n2749_ & new_n2728_;
  assign new_n2753_ = new_n2751_ | new_n2752_;
  assign new_n2754_ = ~new_n2743_;
  assign new_n2755_ = ~new_n2738_;
  assign new_n2756_ = new_n2743_ & new_n2755_;
  assign new_n2757_ = new_n2754_ & new_n2738_;
  assign new_n2758_ = new_n2756_ | new_n2757_;
  assign new_n2759_ = ~new_n2753_;
  assign new_n2760_ = ~new_n2748_;
  assign new_n2761_ = new_n2753_ & new_n2760_;
  assign new_n2762_ = new_n2759_ & new_n2748_;
  assign new_n2763_ = new_n2761_ | new_n2762_;
  assign new_n2764_ = ~pi255;
  assign new_n2765_ = ~new_n2758_;
  assign new_n2766_ = pi255 & new_n2765_;
  assign new_n2767_ = new_n2764_ & new_n2758_;
  assign new_n2768_ = new_n2766_ | new_n2767_;
  assign new_n2769_ = ~pi256;
  assign new_n2770_ = ~new_n2763_;
  assign new_n2771_ = pi256 & new_n2770_;
  assign new_n2772_ = new_n2769_ & new_n2763_;
  assign new_n2773_ = new_n2771_ | new_n2772_;
  assign new_n2774_ = ~po197;
  assign new_n2775_ = ~po198;
  assign new_n2776_ = po197 & new_n2775_;
  assign new_n2777_ = new_n2774_ & po198;
  assign new_n2778_ = new_n2776_ | new_n2777_;
  assign new_n2779_ = ~po195;
  assign new_n2780_ = ~po196;
  assign new_n2781_ = po195 & new_n2780_;
  assign new_n2782_ = new_n2779_ & po196;
  assign new_n2783_ = new_n2781_ | new_n2782_;
  assign new_n2784_ = ~po193;
  assign new_n2785_ = ~po194;
  assign new_n2786_ = po193 & new_n2785_;
  assign new_n2787_ = new_n2784_ & po194;
  assign new_n2788_ = new_n2786_ | new_n2787_;
  assign new_n2789_ = ~po199;
  assign new_n2790_ = ~po206;
  assign new_n2791_ = po199 & new_n2790_;
  assign new_n2792_ = new_n2789_ & po206;
  assign new_n2793_ = new_n2791_ | new_n2792_;
  assign new_n2794_ = ~po204;
  assign new_n2795_ = ~po205;
  assign new_n2796_ = po204 & new_n2795_;
  assign new_n2797_ = new_n2794_ & po205;
  assign new_n2798_ = new_n2796_ | new_n2797_;
  assign new_n2799_ = ~po202;
  assign new_n2800_ = ~po203;
  assign new_n2801_ = po202 & new_n2800_;
  assign new_n2802_ = new_n2799_ & po203;
  assign new_n2803_ = new_n2801_ | new_n2802_;
  assign new_n2804_ = ~po200;
  assign new_n2805_ = ~po201;
  assign new_n2806_ = po200 & new_n2805_;
  assign new_n2807_ = new_n2804_ & po201;
  assign new_n2808_ = new_n2806_ | new_n2807_;
  assign new_n2809_ = ~po207;
  assign new_n2810_ = ~po208;
  assign new_n2811_ = po207 & new_n2810_;
  assign new_n2812_ = new_n2809_ & po208;
  assign new_n2813_ = new_n2811_ | new_n2812_;
  assign new_n2814_ = ~new_n2783_;
  assign new_n2815_ = ~new_n2778_;
  assign new_n2816_ = new_n2783_ & new_n2815_;
  assign new_n2817_ = new_n2814_ & new_n2778_;
  assign new_n2818_ = new_n2816_ | new_n2817_;
  assign new_n2819_ = ~new_n2793_;
  assign new_n2820_ = ~new_n2788_;
  assign new_n2821_ = new_n2793_ & new_n2820_;
  assign new_n2822_ = new_n2819_ & new_n2788_;
  assign new_n2823_ = new_n2821_ | new_n2822_;
  assign new_n2824_ = ~new_n2803_;
  assign new_n2825_ = ~new_n2798_;
  assign new_n2826_ = new_n2803_ & new_n2825_;
  assign new_n2827_ = new_n2824_ & new_n2798_;
  assign new_n2828_ = new_n2826_ | new_n2827_;
  assign new_n2829_ = ~new_n2813_;
  assign new_n2830_ = ~new_n2808_;
  assign new_n2831_ = new_n2813_ & new_n2830_;
  assign new_n2832_ = new_n2829_ & new_n2808_;
  assign new_n2833_ = new_n2831_ | new_n2832_;
  assign new_n2834_ = ~new_n2823_;
  assign new_n2835_ = ~new_n2818_;
  assign new_n2836_ = new_n2823_ & new_n2835_;
  assign new_n2837_ = new_n2834_ & new_n2818_;
  assign new_n2838_ = new_n2836_ | new_n2837_;
  assign new_n2839_ = ~new_n2833_;
  assign new_n2840_ = ~new_n2828_;
  assign new_n2841_ = new_n2833_ & new_n2840_;
  assign new_n2842_ = new_n2839_ & new_n2828_;
  assign new_n2843_ = new_n2841_ | new_n2842_;
  assign new_n2844_ = ~pi128;
  assign new_n2845_ = ~new_n1876_;
  assign new_n2846_ = pi128 & new_n2845_;
  assign new_n2847_ = new_n2844_ & new_n1876_;
  assign new_n2848_ = new_n2846_ | new_n2847_;
  assign new_n2849_ = ~pi127;
  assign new_n2850_ = ~new_n1877_;
  assign new_n2851_ = pi127 & new_n2850_;
  assign new_n2852_ = new_n2849_ & new_n1877_;
  assign new_n2853_ = new_n2851_ | new_n2852_;
  assign new_n2854_ = ~pi126;
  assign new_n2855_ = ~new_n1878_;
  assign new_n2856_ = pi126 & new_n2855_;
  assign new_n2857_ = new_n2854_ & new_n1878_;
  assign new_n2858_ = new_n2856_ | new_n2857_;
  assign new_n2859_ = ~pi125;
  assign new_n2860_ = ~new_n1879_;
  assign new_n2861_ = pi125 & new_n2860_;
  assign new_n2862_ = new_n2859_ & new_n1879_;
  assign new_n2863_ = new_n2861_ | new_n2862_;
  assign new_n2864_ = ~pi124;
  assign new_n2865_ = ~new_n1880_;
  assign new_n2866_ = pi124 & new_n2865_;
  assign new_n2867_ = new_n2864_ & new_n1880_;
  assign new_n2868_ = new_n2866_ | new_n2867_;
  assign new_n2869_ = ~pi123;
  assign new_n2870_ = ~new_n1881_;
  assign new_n2871_ = pi123 & new_n2870_;
  assign new_n2872_ = new_n2869_ & new_n1881_;
  assign new_n2873_ = new_n2871_ | new_n2872_;
  assign new_n2874_ = ~pi122;
  assign new_n2875_ = ~new_n1882_;
  assign new_n2876_ = pi122 & new_n2875_;
  assign new_n2877_ = new_n2874_ & new_n1882_;
  assign new_n2878_ = new_n2876_ | new_n2877_;
  assign new_n2879_ = ~pi121;
  assign new_n2880_ = ~new_n1883_;
  assign new_n2881_ = pi121 & new_n2880_;
  assign new_n2882_ = new_n2879_ & new_n1883_;
  assign new_n2883_ = new_n2881_ | new_n2882_;
  assign new_n2884_ = ~pi120;
  assign new_n2885_ = ~pi119;
  assign new_n2886_ = pi120 & new_n2885_;
  assign new_n2887_ = new_n2884_ & pi119;
  assign new_n2888_ = new_n2886_ | new_n2887_;
  assign new_n2889_ = ~pi011;
  assign new_n2890_ = ~pi010;
  assign new_n2891_ = pi011 & new_n2890_;
  assign new_n2892_ = new_n2889_ & pi010;
  assign new_n2893_ = new_n2891_ | new_n2892_;
  assign new_n2894_ = ~pi109;
  assign new_n2895_ = ~pi110;
  assign new_n2896_ = pi109 & new_n2895_;
  assign new_n2897_ = new_n2894_ & pi110;
  assign new_n2898_ = new_n2896_ | new_n2897_;
  assign new_n2899_ = ~pi243;
  assign new_n2900_ = ~pi244;
  assign new_n2901_ = pi243 & new_n2900_;
  assign new_n2902_ = new_n2899_ & pi244;
  assign new_n2903_ = new_n2901_ | new_n2902_;
  assign new_n2904_ = ~new_n1851_;
  assign new_n2905_ = ~new_n1974_;
  assign new_n2906_ = new_n1851_ & new_n2905_;
  assign new_n2907_ = new_n2904_ & new_n1974_;
  assign new_n2908_ = new_n2906_ | new_n2907_;
  assign new_n2909_ = ~new_n1853_;
  assign new_n2910_ = ~new_n1973_;
  assign new_n2911_ = new_n1853_ & new_n2910_;
  assign new_n2912_ = new_n2909_ & new_n1973_;
  assign new_n2913_ = new_n2911_ | new_n2912_;
  assign new_n2914_ = ~new_n1849_;
  assign new_n2915_ = ~new_n1971_;
  assign new_n2916_ = new_n1849_ & new_n2915_;
  assign new_n2917_ = new_n2914_ & new_n1971_;
  assign new_n2918_ = new_n2916_ | new_n2917_;
  assign new_n2919_ = ~new_n2913_;
  assign new_n2920_ = ~new_n2021_;
  assign new_n2921_ = new_n2913_ & new_n2920_;
  assign new_n2922_ = new_n2919_ & new_n2021_;
  assign new_n2923_ = new_n2921_ | new_n2922_;
  assign new_n2924_ = ~new_n2025_;
  assign new_n2925_ = ~new_n2918_;
  assign new_n2926_ = new_n2025_ & new_n2925_;
  assign new_n2927_ = new_n2924_ & new_n2918_;
  assign new_n2928_ = new_n2926_ | new_n2927_;
  assign new_n2929_ = ~new_n1971_;
  assign new_n2930_ = ~new_n2029_;
  assign new_n2931_ = new_n1971_ & new_n2930_;
  assign new_n2932_ = new_n2929_ & new_n2029_;
  assign new_n2933_ = new_n2931_ | new_n2932_;
  assign new_n2934_ = ~new_n2923_;
  assign new_n2935_ = ~new_n2030_;
  assign new_n2936_ = new_n2923_ & new_n2935_;
  assign new_n2937_ = new_n2934_ & new_n2030_;
  assign new_n2938_ = new_n2936_ | new_n2937_;
  assign new_n2939_ = ~new_n2928_;
  assign new_n2940_ = ~new_n2033_;
  assign new_n2941_ = new_n2928_ & new_n2940_;
  assign new_n2942_ = new_n2939_ & new_n2033_;
  assign new_n2943_ = new_n2941_ | new_n2942_;
  assign new_n2944_ = ~new_n2933_;
  assign new_n2945_ = ~new_n2034_;
  assign new_n2946_ = new_n2933_ & new_n2945_;
  assign new_n2947_ = new_n2944_ & new_n2034_;
  assign new_n2948_ = new_n2946_ | new_n2947_;
  assign new_n2949_ = ~new_n2938_;
  assign new_n2950_ = ~new_n2035_;
  assign new_n2951_ = new_n2938_ & new_n2950_;
  assign new_n2952_ = new_n2949_ & new_n2035_;
  assign new_n2953_ = new_n2951_ | new_n2952_;
  assign new_n2954_ = ~new_n2943_;
  assign new_n2955_ = ~new_n2038_;
  assign new_n2956_ = new_n2943_ & new_n2955_;
  assign new_n2957_ = new_n2954_ & new_n2038_;
  assign new_n2958_ = new_n2956_ | new_n2957_;
  assign new_n2959_ = ~new_n2948_;
  assign new_n2960_ = ~new_n2039_;
  assign new_n2961_ = new_n2948_ & new_n2960_;
  assign new_n2962_ = new_n2959_ & new_n2039_;
  assign new_n2963_ = new_n2961_ | new_n2962_;
  assign new_n2964_ = ~new_n2048_;
  assign new_n2965_ = ~new_n2052_;
  assign new_n2966_ = new_n2048_ & new_n2965_;
  assign new_n2967_ = new_n2964_ & new_n2052_;
  assign new_n2968_ = new_n2966_ | new_n2967_;
  assign new_n2969_ = ~new_n2045_;
  assign new_n2970_ = ~new_n2055_;
  assign new_n2971_ = new_n2045_ & new_n2970_;
  assign new_n2972_ = new_n2969_ & new_n2055_;
  assign new_n2973_ = new_n2971_ | new_n2972_;
  assign new_n2974_ = ~new_n2042_;
  assign new_n2975_ = ~new_n2056_;
  assign new_n2976_ = new_n2042_ & new_n2975_;
  assign new_n2977_ = new_n2974_ & new_n2056_;
  assign new_n2978_ = new_n2976_ | new_n2977_;
endmodule


