// Benchmark "C5315.iscas" written by ABC on Thu Mar 19 13:02:36 2020

module C5315_iscas  ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122;
  wire new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_,
    new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_,
    new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n345_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n384_, new_n385_, new_n386_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n479_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_,
    new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n746_, new_n747_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n970_, new_n971_, new_n972_, new_n973_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_,
    new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_,
    new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_,
    new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_,
    new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_,
    new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_,
    new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1403_, new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_,
    new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_,
    new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_,
    new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_,
    new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_,
    new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_,
    new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_,
    new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_,
    new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_,
    new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_,
    new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_,
    new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_,
    new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_,
    new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_,
    new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_,
    new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_,
    new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_,
    new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_,
    new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_,
    new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_,
    new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_,
    new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_,
    new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_,
    new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_,
    new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_,
    new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_,
    new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_,
    new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_,
    new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_,
    new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_,
    new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_,
    new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_,
    new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_,
    new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_,
    new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_,
    new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_,
    new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_,
    new_n1641_, new_n1642_, new_n1644_, new_n1645_, new_n1646_, new_n1647_,
    new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_,
    new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_,
    new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_,
    new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_,
    new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_,
    new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_,
    new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_,
    new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_,
    new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_,
    new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_,
    new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_,
    new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_,
    new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_,
    new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_,
    new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_,
    new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_,
    new_n1744_, new_n1745_, new_n1746_, new_n1748_, new_n1749_, new_n1750_,
    new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_,
    new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_,
    new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_,
    new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_,
    new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_,
    new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_,
    new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_,
    new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_,
    new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_,
    new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_,
    new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1817_,
    new_n1818_, new_n1819_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1875_, new_n1877_, new_n1878_, new_n1879_, new_n1880_,
    new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_,
    new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_,
    new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_,
    new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_,
    new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_,
    new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_,
    new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_,
    new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_,
    new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_,
    new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_,
    new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_,
    new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_,
    new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_,
    new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_,
    new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_,
    new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_,
    new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_,
    new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_,
    new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_,
    new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_,
    new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_,
    new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_,
    new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2019_, new_n2020_,
    new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_,
    new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_,
    new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_,
    new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2045_,
    new_n2046_, new_n2047_, new_n2048_, new_n2051_, new_n2052_, new_n2053_,
    new_n2054_, new_n2055_, new_n2056_, new_n2058_, new_n2059_, new_n2060_,
    new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_,
    new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2072_,
    new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_,
    new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_,
    new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_,
    new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_,
    new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2102_, new_n2103_,
    new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_,
    new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_,
    new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_,
    new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_,
    new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_,
    new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_,
    new_n2140_, new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_,
    new_n2146_, new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2151_,
    new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_,
    new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_,
    new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_,
    new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_,
    new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_,
    new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_,
    new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2195_,
    new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_,
    new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_,
    new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_,
    new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_,
    new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_,
    new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_,
    new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_,
    new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_,
    new_n2244_, new_n2245_, new_n2246_, new_n2253_, new_n2254_, new_n2258_,
    new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_,
    new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_,
    new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2277_,
    new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_, new_n2283_,
    new_n2284_, new_n2285_, new_n2286_, new_n2288_, new_n2289_, new_n2290_,
    new_n2291_, new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_,
    new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2304_, new_n2309_,
    new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_,
    new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_,
    new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_,
    new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_,
    new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_,
    new_n2354_, new_n2355_, new_n2356_, new_n2358_, new_n2359_, new_n2365_,
    new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_,
    new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_, new_n2377_,
    new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_,
    new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2390_,
    new_n2391_, new_n2393_, new_n2394_, new_n2404_, new_n2405_, new_n2406_,
    new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_,
    new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_,
    new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_,
    new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_,
    new_n2437_, new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_,
    new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_,
    new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_,
    new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_,
    new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_,
    new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_,
    new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_,
    new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_,
    new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_,
    new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_,
    new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_,
    new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_,
    new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_,
    new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_,
    new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_,
    new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_,
    new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_,
    new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_,
    new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_,
    new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_,
    new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_,
    new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_,
    new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_,
    new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_,
    new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_,
    new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_,
    new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2605_, new_n2606_;
  assign new_n302_ = pi176;
  assign new_n303_ = pi176;
  assign new_n304_ = pi176;
  assign new_n305_ = pi176;
  assign new_n306_ = pi176;
  assign new_n307_ = pi175;
  assign new_n308_ = pi175;
  assign new_n309_ = pi175;
  assign new_n310_ = pi175;
  assign new_n311_ = pi175;
  assign new_n312_ = pi174;
  assign new_n313_ = pi174;
  assign new_n314_ = pi173;
  assign new_n315_ = pi173;
  assign new_n316_ = pi172;
  assign new_n317_ = pi172;
  assign new_n318_ = pi171;
  assign new_n319_ = pi171;
  assign new_n320_ = ~pi170;
  assign new_n321_ = ~pi169;
  assign new_n322_ = ~pi168;
  assign new_n323_ = ~pi167;
  assign new_n324_ = ~pi166;
  assign new_n325_ = ~pi165;
  assign po002 = pi164;
  assign new_n327_ = ~pi164;
  assign new_n328_ = ~pi163;
  assign new_n329_ = ~pi162;
  assign new_n330_ = pi162;
  assign new_n331_ = ~pi161;
  assign new_n332_ = pi160;
  assign new_n333_ = pi160;
  assign new_n334_ = pi159;
  assign new_n335_ = pi159;
  assign new_n336_ = pi158;
  assign new_n337_ = pi158;
  assign new_n338_ = pi157;
  assign new_n339_ = pi157;
  assign new_n340_ = ~pi156;
  assign po015 = ~pi155;
  assign po016 = ~pi154;
  assign po014 = ~pi152;
  assign po006 = pi152 & pi155;
  assign new_n345_ = pi151;
  assign po007 = ~pi151;
  assign po009 = ~pi150;
  assign po003 = ~pi150;
  assign po008 = ~pi150;
  assign new_n350_ = pi149;
  assign new_n351_ = pi149;
  assign new_n352_ = pi148;
  assign new_n353_ = pi148;
  assign new_n354_ = pi147;
  assign new_n355_ = pi147;
  assign new_n356_ = pi146;
  assign new_n357_ = pi146;
  assign new_n358_ = pi145;
  assign new_n359_ = pi145;
  assign new_n360_ = pi144;
  assign new_n361_ = pi144;
  assign new_n362_ = pi143;
  assign new_n363_ = pi143;
  assign new_n364_ = pi142;
  assign new_n365_ = pi142;
  assign new_n366_ = pi141;
  assign new_n367_ = pi141;
  assign new_n368_ = pi140;
  assign new_n369_ = pi140;
  assign new_n370_ = pi139;
  assign new_n371_ = pi139;
  assign new_n372_ = pi138;
  assign new_n373_ = pi138;
  assign new_n374_ = pi137;
  assign new_n375_ = pi137;
  assign new_n376_ = pi136;
  assign new_n377_ = pi136;
  assign new_n378_ = pi135 & pi153;
  assign new_n379_ = pi152 & pi153 & pi135 & pi154;
  assign new_n380_ = pi134;
  assign new_n381_ = pi134;
  assign new_n382_ = pi131;
  assign po005 = ~pi130;
  assign new_n384_ = pi129;
  assign new_n385_ = pi129;
  assign new_n386_ = pi129;
  assign po011 = ~pi128;
  assign new_n388_ = pi127;
  assign new_n389_ = pi127;
  assign new_n390_ = pi127;
  assign new_n391_ = pi127;
  assign new_n392_ = pi127;
  assign po004 = ~pi126;
  assign new_n394_ = pi125;
  assign new_n395_ = pi125;
  assign new_n396_ = pi125;
  assign new_n397_ = pi125;
  assign new_n398_ = pi125;
  assign po010 = ~pi124;
  assign new_n400_ = pi123;
  assign new_n401_ = pi123;
  assign new_n402_ = pi122;
  assign new_n403_ = pi122;
  assign new_n404_ = pi120;
  assign new_n405_ = pi120;
  assign new_n406_ = pi120;
  assign new_n407_ = pi120;
  assign new_n408_ = ~pi120;
  assign new_n409_ = pi118;
  assign new_n410_ = pi118;
  assign new_n411_ = pi118;
  assign new_n412_ = pi118;
  assign new_n413_ = pi118;
  assign new_n414_ = pi116;
  assign new_n415_ = pi116;
  assign new_n416_ = pi116;
  assign new_n417_ = pi116;
  assign new_n418_ = pi116;
  assign new_n419_ = pi114;
  assign new_n420_ = pi114;
  assign new_n421_ = pi114;
  assign new_n422_ = pi113;
  assign po001 = pi112;
  assign new_n424_ = pi112;
  assign new_n425_ = pi112;
  assign new_n426_ = pi112;
  assign new_n427_ = pi110;
  assign new_n428_ = pi108;
  assign new_n429_ = pi108;
  assign new_n430_ = pi108;
  assign new_n431_ = pi108;
  assign new_n432_ = pi108;
  assign new_n433_ = pi106;
  assign new_n434_ = pi106;
  assign new_n435_ = pi106;
  assign new_n436_ = pi106;
  assign new_n437_ = pi106;
  assign new_n438_ = pi104;
  assign new_n439_ = pi104;
  assign new_n440_ = pi104;
  assign new_n441_ = pi104;
  assign new_n442_ = pi104;
  assign new_n443_ = pi102;
  assign new_n444_ = pi102;
  assign new_n445_ = pi102;
  assign new_n446_ = pi102;
  assign new_n447_ = pi102;
  assign new_n448_ = pi101;
  assign new_n449_ = pi101;
  assign new_n450_ = pi100;
  assign new_n451_ = pi100;
  assign new_n452_ = pi099;
  assign new_n453_ = pi099;
  assign po013 = ~pi098;
  assign new_n455_ = pi097;
  assign new_n456_ = pi097;
  assign new_n457_ = pi095;
  assign new_n458_ = pi095;
  assign new_n459_ = pi095;
  assign new_n460_ = pi095;
  assign new_n461_ = pi095;
  assign new_n462_ = pi093;
  assign new_n463_ = pi093;
  assign new_n464_ = pi093;
  assign new_n465_ = pi093;
  assign new_n466_ = pi093;
  assign new_n467_ = pi091;
  assign new_n468_ = pi091;
  assign new_n469_ = pi091;
  assign new_n470_ = pi091;
  assign new_n471_ = pi091;
  assign new_n472_ = pi089;
  assign new_n473_ = pi089;
  assign new_n474_ = pi089;
  assign new_n475_ = pi089;
  assign new_n476_ = pi089;
  assign new_n477_ = pi087;
  assign po000 = pi065;
  assign new_n479_ = pi065;
  assign po012 = pi065 & pi066;
  assign new_n481_ = pi063;
  assign new_n482_ = pi063;
  assign new_n483_ = pi061 & pi177;
  assign new_n484_ = pi020;
  assign new_n485_ = pi010 & pi011;
  assign new_n486_ = pi011 & pi010;
  assign new_n487_ = pi001;
  assign new_n488_ = pi000;
  assign new_n489_ = ~pi133 | ~pi000;
  assign new_n490_ = ~new_n302_;
  assign new_n491_ = ~new_n303_;
  assign new_n492_ = new_n309_ & new_n304_;
  assign new_n493_ = ~new_n304_;
  assign new_n494_ = new_n310_ & new_n305_;
  assign new_n495_ = ~new_n305_;
  assign new_n496_ = ~new_n306_;
  assign new_n497_ = ~new_n307_;
  assign new_n498_ = ~new_n308_;
  assign new_n499_ = ~new_n309_;
  assign new_n500_ = ~new_n310_;
  assign new_n501_ = ~new_n311_;
  assign new_n502_ = ~new_n312_;
  assign new_n503_ = ~new_n313_;
  assign new_n504_ = ~new_n314_;
  assign new_n505_ = ~new_n315_;
  assign new_n506_ = ~new_n316_;
  assign new_n507_ = ~new_n317_;
  assign new_n508_ = ~new_n318_;
  assign new_n509_ = ~new_n319_;
  assign new_n510_ = new_n325_ & new_n475_;
  assign new_n511_ = new_n325_ & new_n470_;
  assign new_n512_ = new_n325_ & new_n465_;
  assign new_n513_ = new_n325_ & new_n461_;
  assign new_n514_ = new_n325_ & new_n446_;
  assign new_n515_ = new_n325_ & new_n441_;
  assign new_n516_ = new_n325_ & new_n435_;
  assign new_n517_ = new_n325_ & new_n431_;
  assign new_n518_ = new_n325_ & new_n406_;
  assign new_n519_ = new_n325_ & new_n396_;
  assign new_n520_ = new_n325_ & new_n391_;
  assign new_n521_ = ~new_n329_;
  assign new_n522_ = ~new_n330_;
  assign new_n523_ = ~new_n332_;
  assign new_n524_ = ~new_n333_;
  assign new_n525_ = ~new_n334_;
  assign new_n526_ = ~new_n335_;
  assign new_n527_ = ~new_n336_;
  assign new_n528_ = ~new_n337_;
  assign new_n529_ = ~new_n338_;
  assign new_n530_ = ~new_n339_;
  assign po026 = ~new_n345_;
  assign po024 = new_n345_;
  assign new_n533_ = new_n388_ & new_n453_ & pi149;
  assign new_n534_ = new_n390_ & new_n322_ & pi149;
  assign new_n535_ = ~new_n350_;
  assign new_n536_ = ~new_n351_;
  assign new_n537_ = new_n397_ & new_n322_ & pi148;
  assign new_n538_ = new_n395_ & new_n453_ & pi148;
  assign new_n539_ = ~new_n352_;
  assign new_n540_ = ~new_n353_;
  assign new_n541_ = new_n456_ | pi147;
  assign new_n542_ = new_n453_ & pi147;
  assign new_n543_ = new_n325_ | pi147;
  assign new_n544_ = new_n322_ & pi147;
  assign new_n545_ = ~new_n354_;
  assign new_n546_ = ~new_n355_;
  assign new_n547_ = new_n407_ & new_n322_ & pi146;
  assign new_n548_ = new_n405_ & new_n453_ & pi146;
  assign new_n549_ = ~new_n356_;
  assign new_n550_ = ~new_n357_;
  assign new_n551_ = new_n409_ & new_n453_ & pi145;
  assign new_n552_ = new_n411_ & new_n452_ & pi145;
  assign new_n553_ = ~new_n358_;
  assign new_n554_ = ~new_n359_;
  assign new_n555_ = new_n418_ & new_n452_ & pi144;
  assign new_n556_ = new_n416_ & new_n453_ & pi144;
  assign new_n557_ = ~new_n360_;
  assign new_n558_ = ~new_n361_;
  assign new_n559_ = new_n467_ & new_n452_ & pi143;
  assign new_n560_ = new_n469_ & new_n322_ & pi143;
  assign new_n561_ = ~new_n362_;
  assign new_n562_ = ~new_n363_;
  assign new_n563_ = new_n474_ & new_n452_ & pi142;
  assign new_n564_ = new_n476_ & new_n322_ & pi142;
  assign new_n565_ = ~new_n364_;
  assign new_n566_ = ~new_n365_;
  assign new_n567_ = ~new_n366_;
  assign new_n568_ = ~new_n367_;
  assign new_n569_ = new_n457_ & new_n452_ & pi140;
  assign new_n570_ = new_n460_ & new_n322_ & pi140;
  assign new_n571_ = ~new_n368_;
  assign new_n572_ = ~new_n369_;
  assign new_n573_ = new_n464_ & new_n452_ & pi139;
  assign new_n574_ = new_n466_ & new_n322_ & pi139;
  assign new_n575_ = ~new_n370_;
  assign new_n576_ = ~new_n371_;
  assign new_n577_ = new_n436_ & new_n322_ & pi138;
  assign new_n578_ = new_n434_ & new_n452_ & pi138;
  assign new_n579_ = ~new_n372_;
  assign new_n580_ = ~new_n373_;
  assign new_n581_ = new_n438_ & new_n452_ & pi137;
  assign new_n582_ = new_n440_ & new_n322_ & pi137;
  assign new_n583_ = ~new_n374_;
  assign new_n584_ = ~new_n375_;
  assign new_n585_ = new_n447_ & new_n322_ & pi136;
  assign new_n586_ = new_n445_ & new_n452_ & pi136;
  assign new_n587_ = ~new_n376_;
  assign new_n588_ = ~new_n377_;
  assign po020 = ~new_n378_;
  assign new_n590_ = new_n428_ & new_n452_ & pi134;
  assign new_n591_ = new_n430_ & new_n322_ & pi134;
  assign new_n592_ = ~new_n380_;
  assign new_n593_ = ~new_n381_;
  assign new_n594_ = pi132 & new_n403_;
  assign new_n595_ = ~new_n382_;
  assign new_n596_ = pi130 & new_n403_;
  assign new_n597_ = new_n453_ & new_n384_;
  assign new_n598_ = ~new_n384_;
  assign new_n599_ = new_n453_ & new_n385_;
  assign new_n600_ = ~new_n385_;
  assign new_n601_ = ~new_n386_;
  assign new_n602_ = pi128 & new_n403_;
  assign new_n603_ = ~new_n388_;
  assign new_n604_ = new_n456_ & new_n389_;
  assign new_n605_ = ~new_n389_;
  assign new_n606_ = ~new_n390_;
  assign new_n607_ = ~new_n391_;
  assign new_n608_ = ~new_n392_;
  assign new_n609_ = pi126 & new_n403_;
  assign new_n610_ = new_n456_ & new_n394_;
  assign new_n611_ = ~new_n394_;
  assign new_n612_ = ~new_n395_;
  assign new_n613_ = ~new_n396_;
  assign new_n614_ = ~new_n397_;
  assign new_n615_ = ~new_n398_;
  assign new_n616_ = pi124 & new_n403_;
  assign new_n617_ = ~new_n400_;
  assign new_n618_ = ~new_n401_;
  assign new_n619_ = ~new_n402_;
  assign new_n620_ = ~new_n403_;
  assign new_n621_ = pi121 & new_n402_;
  assign new_n622_ = new_n456_ & new_n404_;
  assign new_n623_ = ~new_n404_;
  assign new_n624_ = ~new_n405_;
  assign new_n625_ = ~new_n406_;
  assign new_n626_ = ~new_n407_;
  assign new_n627_ = new_n408_;
  assign new_n628_ = new_n408_;
  assign new_n629_ = pi119 & new_n402_;
  assign new_n630_ = ~new_n409_;
  assign new_n631_ = new_n456_ & new_n410_;
  assign new_n632_ = ~new_n410_;
  assign new_n633_ = ~new_n411_;
  assign new_n634_ = new_n455_ & new_n412_;
  assign new_n635_ = ~new_n412_;
  assign new_n636_ = ~new_n413_;
  assign new_n637_ = pi117 & new_n402_;
  assign new_n638_ = ~new_n414_;
  assign new_n639_ = new_n456_ & new_n415_;
  assign new_n640_ = ~new_n415_;
  assign new_n641_ = ~new_n416_;
  assign new_n642_ = new_n455_ & new_n417_;
  assign new_n643_ = ~new_n417_;
  assign new_n644_ = ~new_n418_;
  assign new_n645_ = pi115 & new_n402_;
  assign new_n646_ = new_n453_ & new_n419_;
  assign new_n647_ = ~new_n419_;
  assign new_n648_ = ~new_n420_;
  assign new_n649_ = new_n452_ & new_n421_;
  assign new_n650_ = ~new_n421_;
  assign new_n651_ = new_n422_;
  assign po025 = new_n422_;
  assign new_n653_ = pi113 & new_n402_;
  assign new_n654_ = ~new_n424_;
  assign new_n655_ = new_n456_ & new_n425_;
  assign new_n656_ = ~new_n425_;
  assign new_n657_ = new_n455_ & new_n426_;
  assign new_n658_ = ~new_n426_;
  assign new_n659_ = pi111 & new_n401_;
  assign new_n660_ = ~new_n427_;
  assign new_n661_ = pi109 & new_n401_;
  assign new_n662_ = ~new_n428_;
  assign new_n663_ = new_n455_ & new_n429_;
  assign new_n664_ = ~new_n429_;
  assign new_n665_ = ~new_n430_;
  assign new_n666_ = ~new_n431_;
  assign new_n667_ = ~new_n432_;
  assign new_n668_ = pi107 & new_n401_;
  assign new_n669_ = new_n455_ & new_n433_;
  assign new_n670_ = ~new_n433_;
  assign new_n671_ = ~new_n434_;
  assign new_n672_ = ~new_n435_;
  assign new_n673_ = ~new_n436_;
  assign new_n674_ = ~new_n437_;
  assign new_n675_ = pi105 & new_n401_;
  assign new_n676_ = ~new_n438_;
  assign new_n677_ = new_n455_ & new_n439_;
  assign new_n678_ = ~new_n439_;
  assign new_n679_ = ~new_n440_;
  assign new_n680_ = ~new_n441_;
  assign new_n681_ = ~new_n442_;
  assign new_n682_ = pi103 & new_n401_;
  assign new_n683_ = ~new_n443_;
  assign new_n684_ = new_n455_ & new_n444_;
  assign new_n685_ = ~new_n444_;
  assign new_n686_ = ~new_n445_;
  assign new_n687_ = ~new_n446_;
  assign new_n688_ = ~new_n447_;
  assign new_n689_ = new_n455_ & new_n473_;
  assign new_n690_ = new_n455_ & new_n468_;
  assign new_n691_ = new_n455_ & new_n463_;
  assign new_n692_ = new_n455_ & new_n458_;
  assign new_n693_ = pi096 & new_n400_;
  assign new_n694_ = ~new_n457_;
  assign new_n695_ = ~new_n458_;
  assign new_n696_ = ~new_n459_;
  assign new_n697_ = ~new_n460_;
  assign new_n698_ = ~new_n461_;
  assign new_n699_ = pi094 & new_n400_;
  assign new_n700_ = ~new_n462_;
  assign new_n701_ = ~new_n463_;
  assign new_n702_ = ~new_n464_;
  assign new_n703_ = ~new_n465_;
  assign new_n704_ = ~new_n466_;
  assign new_n705_ = pi092 & new_n400_;
  assign new_n706_ = ~new_n467_;
  assign new_n707_ = ~new_n468_;
  assign new_n708_ = ~new_n469_;
  assign new_n709_ = ~new_n470_;
  assign new_n710_ = ~new_n471_;
  assign new_n711_ = pi090 & new_n400_;
  assign new_n712_ = ~new_n472_;
  assign new_n713_ = ~new_n473_;
  assign new_n714_ = ~new_n474_;
  assign new_n715_ = ~new_n475_;
  assign new_n716_ = ~new_n476_;
  assign new_n717_ = pi088 & new_n400_;
  assign new_n718_ = new_n477_;
  assign new_n719_ = new_n477_;
  assign new_n720_ = new_n477_;
  assign new_n721_ = new_n477_;
  assign new_n722_ = new_n477_;
  assign new_n723_ = new_n336_ & pi080 & new_n338_;
  assign new_n724_ = new_n332_ & pi080 & new_n334_;
  assign new_n725_ = new_n336_ & pi078 & new_n338_;
  assign new_n726_ = new_n332_ & pi078 & new_n334_;
  assign new_n727_ = new_n333_ & pi076 & new_n335_;
  assign new_n728_ = new_n337_ & pi076 & new_n339_;
  assign new_n729_ = new_n337_ & pi075 & new_n339_;
  assign new_n730_ = new_n333_ & pi075 & new_n335_;
  assign new_n731_ = new_n337_ & pi074 & new_n339_;
  assign new_n732_ = new_n333_ & pi074 & new_n335_;
  assign new_n733_ = new_n333_ & pi073 & new_n335_;
  assign new_n734_ = new_n337_ & pi073 & new_n339_;
  assign new_n735_ = new_n337_ & pi072 & new_n339_;
  assign new_n736_ = new_n333_ & pi072 & new_n335_;
  assign new_n737_ = new_n332_ & pi071 & new_n334_;
  assign new_n738_ = new_n336_ & pi071 & new_n338_;
  assign new_n739_ = new_n336_ & pi069 & new_n338_;
  assign new_n740_ = new_n332_ & pi069 & new_n334_;
  assign new_n741_ = new_n332_ & pi067 & new_n334_;
  assign new_n742_ = new_n336_ & pi067 & new_n338_;
  assign po022 = new_n479_;
  assign new_n744_ = new_n479_;
  assign po027 = ~new_n485_ | ~pi064;
  assign new_n746_ = new_n481_;
  assign new_n747_ = new_n481_;
  assign po021 = new_n481_;
  assign new_n749_ = new_n482_;
  assign new_n750_ = new_n482_;
  assign po018 = pi062 & new_n327_;
  assign new_n752_ = ~new_n483_;
  assign new_n753_ = pi169 & pi053 & new_n320_;
  assign new_n754_ = new_n312_ & pi040 & new_n314_;
  assign new_n755_ = new_n318_ & pi040 & new_n316_;
  assign new_n756_ = new_n312_ & pi039 & new_n314_;
  assign new_n757_ = new_n318_ & pi039 & new_n316_;
  assign new_n758_ = pi037 & new_n306_;
  assign new_n759_ = pi037 & new_n306_;
  assign new_n760_ = pi036 & new_n306_;
  assign new_n761_ = pi036 & new_n306_;
  assign new_n762_ = pi034 & new_n329_;
  assign new_n763_ = pi034 & new_n329_;
  assign new_n764_ = pi032 & new_n329_;
  assign new_n765_ = pi031 & new_n329_;
  assign new_n766_ = new_n313_ & pi024 & new_n315_;
  assign new_n767_ = new_n319_ & pi024 & new_n317_;
  assign new_n768_ = new_n319_ & pi022 & new_n317_;
  assign new_n769_ = new_n313_ & pi022 & new_n315_;
  assign new_n770_ = new_n319_ & pi021 & new_n317_;
  assign new_n771_ = new_n313_ & pi021 & new_n315_;
  assign new_n772_ = ~new_n484_;
  assign new_n773_ = new_n312_ & pi017 & new_n314_;
  assign new_n774_ = new_n318_ & pi017 & new_n316_;
  assign new_n775_ = new_n318_ & pi014 & new_n316_;
  assign new_n776_ = new_n312_ & pi014 & new_n314_;
  assign new_n777_ = new_n312_ & pi013 & new_n314_;
  assign new_n778_ = new_n318_ & pi013 & new_n316_;
  assign po028 = ~new_n485_;
  assign new_n780_ = ~new_n485_;
  assign new_n781_ = new_n328_ & pi010;
  assign new_n782_ = new_n313_ & pi005 & new_n315_;
  assign new_n783_ = new_n319_ & pi005 & new_n317_;
  assign new_n784_ = new_n319_ & pi004 & new_n317_;
  assign new_n785_ = new_n313_ & pi004 & new_n315_;
  assign new_n786_ = ~new_n487_;
  assign new_n787_ = new_n488_;
  assign po023 = new_n488_;
  assign po017 = ~new_n489_;
  assign new_n790_ = new_n324_ & new_n715_;
  assign new_n791_ = new_n324_ & new_n709_;
  assign new_n792_ = new_n324_ & new_n703_;
  assign new_n793_ = new_n324_ & new_n698_;
  assign new_n794_ = new_n324_ & new_n687_;
  assign new_n795_ = new_n324_ & new_n680_;
  assign new_n796_ = new_n324_ & new_n672_;
  assign new_n797_ = new_n324_ & new_n666_;
  assign new_n798_ = new_n324_ & new_n625_;
  assign new_n799_ = new_n324_ & new_n613_;
  assign new_n800_ = new_n324_ & new_n607_;
  assign new_n801_ = new_n330_ & new_n780_;
  assign new_n802_ = new_n330_ & new_n780_;
  assign new_n803_ = new_n330_ & new_n780_;
  assign new_n804_ = new_n330_ & new_n780_;
  assign new_n805_ = new_n522_ & new_n780_;
  assign new_n806_ = new_n522_ & new_n780_;
  assign new_n807_ = new_n522_ & new_n780_;
  assign new_n808_ = new_n522_ & new_n780_;
  assign new_n809_ = new_n603_ & pi149 & new_n451_;
  assign new_n810_ = new_n606_ & pi149 & new_n323_;
  assign new_n811_ = new_n614_ & pi148 & new_n323_;
  assign new_n812_ = new_n612_ & pi148 & new_n451_;
  assign new_n813_ = ~new_n542_;
  assign new_n814_ = ~new_n544_;
  assign new_n815_ = new_n626_ & pi146 & new_n323_;
  assign new_n816_ = new_n624_ & pi146 & new_n451_;
  assign new_n817_ = new_n630_ & pi145 & new_n451_;
  assign new_n818_ = new_n633_ & pi145 & new_n450_;
  assign new_n819_ = new_n644_ & pi144 & new_n450_;
  assign new_n820_ = new_n641_ & pi144 & new_n451_;
  assign new_n821_ = new_n706_ & pi143 & new_n450_;
  assign new_n822_ = new_n708_ & pi143 & new_n323_;
  assign new_n823_ = new_n714_ & pi142 & new_n450_;
  assign new_n824_ = new_n716_ & pi142 & new_n323_;
  assign new_n825_ = new_n721_ & new_n453_ & pi141;
  assign new_n826_ = new_n719_ & new_n453_ & pi141;
  assign new_n827_ = new_n694_ & pi140 & new_n450_;
  assign new_n828_ = new_n697_ & pi140 & new_n323_;
  assign new_n829_ = new_n702_ & pi139 & new_n450_;
  assign new_n830_ = new_n704_ & pi139 & new_n323_;
  assign new_n831_ = new_n673_ & pi138 & new_n323_;
  assign new_n832_ = new_n671_ & pi138 & new_n450_;
  assign new_n833_ = new_n676_ & pi137 & new_n450_;
  assign new_n834_ = new_n679_ & pi137 & new_n323_;
  assign new_n835_ = new_n688_ & pi136 & new_n323_;
  assign new_n836_ = new_n686_ & pi136 & new_n450_;
  assign new_n837_ = new_n662_ & pi134 & new_n450_;
  assign new_n838_ = new_n665_ & pi134 & new_n323_;
  assign new_n839_ = pi131 & new_n620_;
  assign new_n840_ = ~new_n382_ | ~new_n601_;
  assign new_n841_ = pi129 & new_n620_;
  assign new_n842_ = ~new_n386_ | ~new_n595_;
  assign new_n843_ = pi127 & new_n620_;
  assign new_n844_ = ~new_n392_ | ~new_n615_;
  assign new_n845_ = pi125 & new_n620_;
  assign new_n846_ = ~new_n398_ | ~new_n608_;
  assign new_n847_ = new_n620_ | new_n616_;
  assign new_n848_ = pi120 & new_n619_;
  assign new_n849_ = ~new_n627_;
  assign new_n850_ = ~new_n628_;
  assign new_n851_ = pi118 & new_n619_;
  assign new_n852_ = ~new_n413_ | ~new_n638_;
  assign new_n853_ = ~new_n414_ | ~new_n636_;
  assign new_n854_ = pi116 & new_n619_;
  assign new_n855_ = ~new_n420_ | ~new_n654_;
  assign new_n856_ = pi114 & new_n619_;
  assign po034 = ~new_n651_;
  assign po033 = new_n651_;
  assign new_n859_ = ~new_n424_ | ~new_n648_;
  assign new_n860_ = pi112 & new_n619_;
  assign new_n861_ = pi110 & new_n618_;
  assign new_n862_ = ~new_n427_ | ~new_n667_;
  assign new_n863_ = pi108 & new_n618_;
  assign new_n864_ = ~new_n432_ | ~new_n660_;
  assign new_n865_ = pi106 & new_n618_;
  assign new_n866_ = ~new_n437_ | ~new_n681_;
  assign new_n867_ = pi104 & new_n618_;
  assign new_n868_ = ~new_n442_ | ~new_n674_;
  assign new_n869_ = ~new_n443_ | ~new_n696_;
  assign new_n870_ = pi102 & new_n618_;
  assign new_n871_ = new_n448_ & new_n658_;
  assign new_n872_ = new_n448_ & new_n643_;
  assign new_n873_ = new_n448_ & new_n635_;
  assign new_n874_ = new_n448_ & new_n685_;
  assign new_n875_ = new_n448_ & new_n678_;
  assign new_n876_ = new_n448_ & new_n670_;
  assign new_n877_ = new_n448_ & new_n664_;
  assign new_n878_ = new_n448_ & new_n713_;
  assign new_n879_ = new_n448_ & new_n707_;
  assign new_n880_ = new_n448_ & new_n701_;
  assign new_n881_ = new_n448_ & new_n695_;
  assign new_n882_ = new_n449_ & new_n623_;
  assign new_n883_ = new_n449_ & new_n605_;
  assign new_n884_ = new_n449_ & new_n611_;
  assign new_n885_ = new_n449_ & new_n656_;
  assign new_n886_ = new_n449_ & new_n632_;
  assign new_n887_ = new_n449_ & new_n640_;
  assign new_n888_ = new_n450_ & new_n650_;
  assign new_n889_ = new_n451_ & new_n598_;
  assign new_n890_ = new_n451_ & new_n600_;
  assign new_n891_ = new_n451_ & new_n647_;
  assign new_n892_ = new_n456_ & new_n718_;
  assign new_n893_ = new_n456_ & new_n720_;
  assign new_n894_ = pi095 & new_n617_;
  assign new_n895_ = ~new_n459_ | ~new_n683_;
  assign new_n896_ = ~new_n462_ | ~new_n710_;
  assign new_n897_ = pi093 & new_n617_;
  assign new_n898_ = pi091 & new_n617_;
  assign new_n899_ = ~new_n471_ | ~new_n700_;
  assign new_n900_ = ~new_n722_ | ~new_n712_;
  assign new_n901_ = pi089 & new_n617_;
  assign new_n902_ = ~new_n718_;
  assign new_n903_ = ~new_n719_;
  assign new_n904_ = ~new_n720_;
  assign new_n905_ = ~new_n721_;
  assign new_n906_ = ~new_n722_;
  assign new_n907_ = pi087 & new_n617_;
  assign new_n908_ = new_n333_ & pi086 & new_n526_;
  assign new_n909_ = new_n337_ & pi086 & new_n530_;
  assign new_n910_ = new_n333_ & pi085 & new_n526_;
  assign new_n911_ = new_n337_ & pi085 & new_n530_;
  assign new_n912_ = new_n333_ & pi084 & new_n526_;
  assign new_n913_ = new_n337_ & pi084 & new_n530_;
  assign new_n914_ = new_n333_ & pi083 & new_n526_;
  assign new_n915_ = new_n337_ & pi083 & new_n530_;
  assign new_n916_ = new_n333_ & pi082 & new_n526_;
  assign new_n917_ = new_n337_ & pi082 & new_n530_;
  assign new_n918_ = new_n336_ & pi081 & new_n529_;
  assign new_n919_ = new_n332_ & pi081 & new_n525_;
  assign new_n920_ = new_n332_ & pi079 & new_n525_;
  assign new_n921_ = new_n336_ & pi079 & new_n529_;
  assign new_n922_ = new_n332_ & pi077 & new_n525_;
  assign new_n923_ = new_n336_ & pi077 & new_n529_;
  assign new_n924_ = new_n332_ & pi070 & new_n525_;
  assign new_n925_ = new_n336_ & pi070 & new_n529_;
  assign new_n926_ = new_n336_ & pi068 & new_n529_;
  assign new_n927_ = new_n332_ & pi068 & new_n525_;
  assign new_n928_ = new_n304_ & pi059 & new_n499_;
  assign new_n929_ = new_n304_ & pi058 & new_n499_;
  assign new_n930_ = new_n304_ & pi057 & new_n499_;
  assign new_n931_ = new_n305_ & pi056 & new_n500_;
  assign new_n932_ = new_n305_ & pi055 & new_n500_;
  assign new_n933_ = new_n305_ & pi054 & new_n500_;
  assign new_n934_ = new_n302_ & pi053 & new_n497_;
  assign new_n935_ = new_n303_ & pi052 & new_n498_;
  assign new_n936_ = new_n302_ & pi051 & new_n497_;
  assign new_n937_ = new_n304_ & pi050 & new_n499_;
  assign new_n938_ = new_n304_ & pi049 & new_n499_;
  assign new_n939_ = new_n305_ & pi048 & new_n500_;
  assign new_n940_ = new_n305_ & pi047 & new_n500_;
  assign new_n941_ = new_n302_ & pi046 & new_n497_;
  assign new_n942_ = new_n303_ & pi045 & new_n498_;
  assign new_n943_ = new_n303_ & pi044 & new_n498_;
  assign new_n944_ = new_n303_ & pi043 & new_n498_;
  assign new_n945_ = new_n302_ & pi042 & new_n497_;
  assign new_n946_ = new_n312_ & pi041 & new_n504_;
  assign new_n947_ = new_n318_ & pi041 & new_n506_;
  assign new_n948_ = new_n312_ & pi038 & new_n504_;
  assign new_n949_ = new_n318_ & pi038 & new_n506_;
  assign new_n950_ = new_n312_ & pi035 & new_n504_;
  assign new_n951_ = new_n318_ & pi035 & new_n506_;
  assign new_n952_ = pi033 & new_n521_;
  assign new_n953_ = pi031 & new_n521_;
  assign new_n954_ = new_n313_ & pi026 & new_n505_;
  assign new_n955_ = new_n319_ & pi026 & new_n507_;
  assign new_n956_ = new_n319_ & pi025 & new_n507_;
  assign new_n957_ = new_n313_ & pi025 & new_n505_;
  assign new_n958_ = new_n313_ & pi023 & new_n505_;
  assign new_n959_ = new_n319_ & pi023 & new_n507_;
  assign new_n960_ = new_n303_ & pi019 & new_n498_;
  assign new_n961_ = new_n302_ & pi018 & new_n497_;
  assign new_n962_ = new_n312_ & pi016 & new_n504_;
  assign new_n963_ = new_n318_ & pi016 & new_n506_;
  assign new_n964_ = new_n312_ & pi015 & new_n504_;
  assign new_n965_ = new_n318_ & pi015 & new_n506_;
  assign new_n966_ = pi012 & new_n521_;
  assign new_n967_ = pi012 & new_n521_;
  assign new_n968_ = ~new_n780_;
  assign po019 = ~new_n781_;
  assign new_n970_ = new_n313_ & pi003 & new_n505_;
  assign new_n971_ = new_n319_ & pi003 & new_n507_;
  assign new_n972_ = new_n319_ & pi002 & new_n507_;
  assign new_n973_ = new_n313_ & pi002 & new_n505_;
  assign po029 = new_n787_;
  assign po030 = new_n787_;
  assign po031 = new_n787_;
  assign po032 = new_n787_;
  assign new_n978_ = pi149 | new_n604_ | new_n883_;
  assign new_n979_ = new_n533_ | new_n809_;
  assign new_n980_ = pi149 | new_n520_ | new_n800_;
  assign new_n981_ = new_n534_ | new_n810_;
  assign new_n982_ = new_n537_ | new_n811_;
  assign new_n983_ = pi148 | new_n519_ | new_n799_;
  assign new_n984_ = new_n538_ | new_n812_;
  assign new_n985_ = pi148 | new_n610_ | new_n884_;
  assign new_n986_ = new_n813_ & new_n541_;
  assign new_n987_ = new_n814_ & new_n543_;
  assign new_n988_ = pi147 & new_n847_;
  assign new_n989_ = new_n847_ & pi147;
  assign new_n990_ = new_n547_ | new_n815_;
  assign new_n991_ = pi146 | new_n518_ | new_n798_;
  assign new_n992_ = new_n548_ | new_n816_;
  assign new_n993_ = pi146 | new_n622_ | new_n882_;
  assign new_n994_ = pi145 | new_n631_ | new_n886_;
  assign new_n995_ = new_n551_ | new_n817_;
  assign new_n996_ = pi145 | new_n634_ | new_n873_;
  assign new_n997_ = new_n552_ | new_n818_;
  assign new_n998_ = new_n555_ | new_n819_;
  assign new_n999_ = pi144 | new_n642_ | new_n872_;
  assign new_n1000_ = new_n556_ | new_n820_;
  assign new_n1001_ = pi144 | new_n639_ | new_n887_;
  assign new_n1002_ = pi143 | new_n690_ | new_n879_;
  assign new_n1003_ = new_n559_ | new_n821_;
  assign new_n1004_ = pi143 | new_n511_ | new_n791_;
  assign new_n1005_ = new_n560_ | new_n822_;
  assign new_n1006_ = new_n563_ | new_n823_;
  assign new_n1007_ = pi142 | new_n689_ | new_n878_;
  assign new_n1008_ = new_n564_ | new_n824_;
  assign new_n1009_ = pi142 | new_n510_ | new_n790_;
  assign new_n1010_ = new_n905_ & pi141 & new_n451_;
  assign new_n1011_ = new_n903_ & pi141 & new_n451_;
  assign new_n1012_ = pi140 | new_n692_ | new_n881_;
  assign new_n1013_ = new_n569_ | new_n827_;
  assign new_n1014_ = pi140 | new_n513_ | new_n793_;
  assign new_n1015_ = new_n570_ | new_n828_;
  assign new_n1016_ = new_n573_ | new_n829_;
  assign new_n1017_ = pi139 | new_n691_ | new_n880_;
  assign new_n1018_ = new_n574_ | new_n830_;
  assign new_n1019_ = pi139 | new_n512_ | new_n792_;
  assign new_n1020_ = new_n577_ | new_n831_;
  assign new_n1021_ = pi138 | new_n516_ | new_n796_;
  assign new_n1022_ = new_n578_ | new_n832_;
  assign new_n1023_ = pi138 | new_n669_ | new_n876_;
  assign new_n1024_ = pi137 | new_n677_ | new_n875_;
  assign new_n1025_ = new_n581_ | new_n833_;
  assign new_n1026_ = pi137 | new_n515_ | new_n795_;
  assign new_n1027_ = new_n582_ | new_n834_;
  assign new_n1028_ = new_n585_ | new_n835_;
  assign new_n1029_ = pi136 | new_n514_ | new_n794_;
  assign new_n1030_ = new_n586_ | new_n836_;
  assign new_n1031_ = pi136 | new_n684_ | new_n874_;
  assign new_n1032_ = pi134 | new_n663_ | new_n877_;
  assign new_n1033_ = new_n590_ | new_n837_;
  assign new_n1034_ = pi134 | new_n517_ | new_n797_;
  assign new_n1035_ = new_n591_ | new_n838_;
  assign new_n1036_ = new_n839_ | new_n594_;
  assign new_n1037_ = ~new_n840_ | ~new_n842_;
  assign new_n1038_ = new_n841_ | new_n596_;
  assign new_n1039_ = new_n597_ | new_n889_;
  assign new_n1040_ = new_n599_ | new_n890_;
  assign new_n1041_ = new_n843_ | new_n602_;
  assign new_n1042_ = ~new_n844_ | ~new_n846_;
  assign new_n1043_ = new_n845_ | new_n609_;
  assign new_n1044_ = new_n847_;
  assign new_n1045_ = new_n847_;
  assign new_n1046_ = new_n847_;
  assign new_n1047_ = new_n848_ | new_n621_;
  assign new_n1048_ = new_n851_ | new_n629_;
  assign new_n1049_ = ~new_n852_ | ~new_n853_;
  assign new_n1050_ = new_n854_ | new_n637_;
  assign new_n1051_ = new_n856_ | new_n645_;
  assign new_n1052_ = new_n646_ | new_n891_;
  assign new_n1053_ = ~new_n855_ | ~new_n859_;
  assign new_n1054_ = new_n649_ | new_n888_;
  assign new_n1055_ = new_n860_ | new_n653_;
  assign new_n1056_ = new_n655_ | new_n885_;
  assign new_n1057_ = new_n657_ | new_n871_;
  assign new_n1058_ = new_n861_ | new_n659_;
  assign new_n1059_ = ~new_n862_ | ~new_n864_;
  assign new_n1060_ = new_n863_ | new_n661_;
  assign new_n1061_ = new_n865_ | new_n668_;
  assign new_n1062_ = ~new_n866_ | ~new_n868_;
  assign new_n1063_ = new_n867_ | new_n675_;
  assign new_n1064_ = new_n870_ | new_n682_;
  assign new_n1065_ = ~new_n869_ | ~new_n895_;
  assign new_n1066_ = new_n449_ & new_n902_;
  assign new_n1067_ = new_n449_ & new_n904_;
  assign new_n1068_ = new_n894_ | new_n693_;
  assign new_n1069_ = new_n897_ | new_n699_;
  assign new_n1070_ = ~new_n896_ | ~new_n899_;
  assign new_n1071_ = new_n898_ | new_n705_;
  assign new_n1072_ = new_n901_ | new_n711_;
  assign new_n1073_ = ~new_n472_ | ~new_n906_;
  assign new_n1074_ = new_n907_ | new_n717_;
  assign new_n1075_ = new_n966_ | new_n762_;
  assign new_n1076_ = new_n967_ | new_n763_;
  assign new_n1077_ = new_n952_ | new_n764_;
  assign new_n1078_ = new_n953_ | new_n765_;
  assign new_n1079_ = new_n968_ & pi030 & new_n522_;
  assign new_n1080_ = new_n968_ & pi029 & new_n330_;
  assign new_n1081_ = new_n968_ & pi028 & new_n330_;
  assign new_n1082_ = new_n968_ & pi027 & new_n522_;
  assign new_n1083_ = new_n968_ & pi009 & new_n522_;
  assign new_n1084_ = new_n968_ & pi008 & new_n330_;
  assign new_n1085_ = new_n968_ & pi007 & new_n522_;
  assign new_n1086_ = new_n968_ & pi006 & new_n330_;
  assign new_n1087_ = new_n493_ & new_n987_ & new_n499_;
  assign new_n1088_ = new_n801_ | new_n805_ | new_n1082_ | new_n1086_;
  assign new_n1089_ = new_n802_ | new_n808_ | new_n1085_ | new_n1084_;
  assign new_n1090_ = new_n803_ | new_n807_ | new_n1083_ | new_n1080_;
  assign new_n1091_ = new_n804_ | new_n806_ | new_n1079_ | new_n1081_;
  assign new_n1092_ = ~new_n979_;
  assign new_n1093_ = ~new_n981_;
  assign new_n1094_ = pi149 & new_n1041_;
  assign new_n1095_ = new_n1041_ & pi149;
  assign new_n1096_ = ~new_n982_;
  assign new_n1097_ = ~new_n984_;
  assign new_n1098_ = new_n1043_ & pi148;
  assign new_n1099_ = pi148 & new_n1043_;
  assign new_n1100_ = ~new_n986_;
  assign new_n1101_ = ~new_n987_;
  assign new_n1102_ = ~new_n1045_ | ~new_n545_;
  assign new_n1103_ = ~new_n1044_ | ~new_n546_;
  assign new_n1104_ = ~new_n990_;
  assign new_n1105_ = ~new_n992_;
  assign new_n1106_ = pi146 & new_n1047_;
  assign new_n1107_ = new_n1047_ & pi146;
  assign new_n1108_ = ~new_n995_;
  assign new_n1109_ = ~new_n997_;
  assign new_n1110_ = ~pi145 & ~new_n1048_;
  assign new_n1111_ = pi145 & new_n1048_;
  assign new_n1112_ = pi145 & new_n1048_;
  assign new_n1113_ = ~pi145 & ~new_n1048_;
  assign new_n1114_ = ~new_n998_;
  assign new_n1115_ = ~new_n1000_;
  assign new_n1116_ = new_n1050_ & pi144;
  assign new_n1117_ = pi144 & new_n1050_;
  assign new_n1118_ = ~new_n1003_;
  assign new_n1119_ = ~new_n1005_;
  assign new_n1120_ = new_n1071_ & pi143;
  assign new_n1121_ = pi143 & new_n1071_;
  assign new_n1122_ = ~new_n1006_;
  assign new_n1123_ = ~new_n1008_;
  assign new_n1124_ = pi142 & new_n1072_;
  assign new_n1125_ = new_n1072_ & pi142;
  assign new_n1126_ = pi141 | new_n893_ | new_n1067_;
  assign new_n1127_ = new_n825_ | new_n1010_;
  assign new_n1128_ = pi141 | new_n892_ | new_n1066_;
  assign new_n1129_ = new_n826_ | new_n1011_;
  assign new_n1130_ = new_n1074_ & pi141;
  assign new_n1131_ = pi141 & new_n1074_;
  assign new_n1132_ = ~new_n1013_;
  assign new_n1133_ = ~new_n1015_;
  assign new_n1134_ = pi140 & new_n1068_;
  assign new_n1135_ = new_n1068_ & pi140;
  assign new_n1136_ = ~new_n1016_;
  assign new_n1137_ = ~new_n1018_;
  assign new_n1138_ = pi139 & new_n1069_;
  assign new_n1139_ = ~pi139 & ~new_n1069_;
  assign new_n1140_ = ~pi139 & ~new_n1069_;
  assign new_n1141_ = pi139 & new_n1069_;
  assign new_n1142_ = ~new_n1020_;
  assign new_n1143_ = ~new_n1022_;
  assign new_n1144_ = new_n1061_ & pi138;
  assign new_n1145_ = pi138 & new_n1061_;
  assign new_n1146_ = ~new_n1025_;
  assign new_n1147_ = ~new_n1027_;
  assign new_n1148_ = pi137 & new_n1063_;
  assign new_n1149_ = new_n1063_ & pi137;
  assign new_n1150_ = ~new_n1028_;
  assign new_n1151_ = ~new_n1030_;
  assign new_n1152_ = new_n1064_ & pi136;
  assign new_n1153_ = pi136 & new_n1064_;
  assign new_n1154_ = ~new_n1033_;
  assign new_n1155_ = ~new_n1035_;
  assign new_n1156_ = ~pi134 & ~new_n1060_;
  assign new_n1157_ = pi134 & new_n1060_;
  assign new_n1158_ = new_n1060_ & pi134;
  assign new_n1159_ = ~new_n1036_;
  assign new_n1160_ = ~new_n1037_;
  assign new_n1161_ = ~new_n1038_;
  assign new_n1162_ = new_n1038_;
  assign new_n1163_ = new_n1038_;
  assign new_n1164_ = ~new_n1038_;
  assign new_n1165_ = new_n1038_;
  assign new_n1166_ = ~new_n1039_;
  assign new_n1167_ = ~new_n1040_;
  assign new_n1168_ = new_n1041_;
  assign new_n1169_ = new_n1041_;
  assign new_n1170_ = new_n1041_;
  assign new_n1171_ = ~new_n1042_;
  assign new_n1172_ = new_n1043_;
  assign new_n1173_ = new_n1043_;
  assign new_n1174_ = new_n1043_;
  assign new_n1175_ = ~new_n1044_;
  assign new_n1176_ = ~new_n1045_;
  assign new_n1177_ = ~new_n1046_;
  assign new_n1178_ = new_n1047_;
  assign new_n1179_ = new_n1047_;
  assign new_n1180_ = new_n1047_;
  assign new_n1181_ = new_n628_ & new_n1042_ & new_n1037_;
  assign new_n1182_ = new_n1048_;
  assign new_n1183_ = new_n1048_;
  assign new_n1184_ = new_n1048_;
  assign new_n1185_ = ~new_n1049_;
  assign new_n1186_ = new_n1050_;
  assign new_n1187_ = new_n1050_;
  assign new_n1188_ = new_n1050_;
  assign new_n1189_ = ~new_n1051_;
  assign new_n1190_ = new_n1051_;
  assign new_n1191_ = ~new_n1051_;
  assign new_n1192_ = new_n1051_;
  assign new_n1193_ = new_n1051_;
  assign new_n1194_ = ~new_n1052_;
  assign new_n1195_ = ~new_n1053_;
  assign new_n1196_ = ~new_n1054_;
  assign new_n1197_ = ~new_n1055_;
  assign new_n1198_ = ~new_n1055_;
  assign new_n1199_ = new_n1055_;
  assign new_n1200_ = new_n1055_;
  assign new_n1201_ = ~new_n1056_;
  assign new_n1202_ = ~new_n1057_;
  assign new_n1203_ = new_n1057_;
  assign new_n1204_ = ~new_n1058_;
  assign new_n1205_ = ~new_n1059_;
  assign new_n1206_ = new_n1060_;
  assign new_n1207_ = new_n1060_;
  assign new_n1208_ = new_n1060_;
  assign new_n1209_ = new_n1061_;
  assign new_n1210_ = new_n1061_;
  assign new_n1211_ = new_n1061_;
  assign new_n1212_ = ~new_n1062_;
  assign new_n1213_ = new_n1063_;
  assign new_n1214_ = new_n1063_;
  assign new_n1215_ = new_n1063_;
  assign new_n1216_ = new_n1064_;
  assign new_n1217_ = new_n1064_;
  assign new_n1218_ = new_n1064_;
  assign new_n1219_ = new_n1065_;
  assign new_n1220_ = new_n1065_;
  assign new_n1221_ = new_n1068_;
  assign new_n1222_ = new_n1068_;
  assign new_n1223_ = new_n1068_;
  assign new_n1224_ = new_n1069_;
  assign new_n1225_ = new_n1069_;
  assign new_n1226_ = new_n1069_;
  assign new_n1227_ = ~new_n1070_;
  assign new_n1228_ = new_n1071_;
  assign new_n1229_ = new_n1071_;
  assign new_n1230_ = new_n1071_;
  assign new_n1231_ = new_n1072_;
  assign new_n1232_ = new_n1072_;
  assign new_n1233_ = new_n1072_;
  assign new_n1234_ = ~new_n1073_ | ~new_n900_;
  assign new_n1235_ = new_n1074_;
  assign new_n1236_ = new_n1074_;
  assign new_n1237_ = new_n1074_;
  assign new_n1238_ = new_n1077_ & new_n486_;
  assign new_n1239_ = new_n1076_ & new_n486_;
  assign new_n1240_ = new_n1075_ & new_n486_;
  assign new_n1241_ = new_n1078_ & new_n486_;
  assign new_n1242_ = new_n490_ & new_n1196_ & new_n497_;
  assign new_n1243_ = new_n490_ & new_n1203_ & new_n497_;
  assign new_n1244_ = new_n493_ & new_n1166_ & new_n499_;
  assign new_n1245_ = new_n321_ & new_n1203_ & new_n320_;
  assign new_n1246_ = new_n1092_ & new_n978_;
  assign new_n1247_ = new_n1093_ & new_n980_;
  assign new_n1248_ = ~new_n1169_ | ~new_n535_;
  assign new_n1249_ = ~new_n1168_ | ~new_n536_;
  assign new_n1250_ = new_n1096_ & new_n983_;
  assign new_n1251_ = new_n1097_ & new_n985_;
  assign new_n1252_ = ~new_n1174_ | ~new_n539_;
  assign new_n1253_ = ~new_n1173_ | ~new_n540_;
  assign new_n1254_ = ~new_n354_ | ~new_n1176_;
  assign new_n1255_ = ~new_n355_ | ~new_n1175_;
  assign new_n1256_ = new_n1104_ & new_n991_;
  assign new_n1257_ = new_n1105_ & new_n993_;
  assign new_n1258_ = ~new_n1180_ | ~new_n549_;
  assign new_n1259_ = ~new_n1179_ | ~new_n550_;
  assign new_n1260_ = new_n1108_ & new_n994_;
  assign new_n1261_ = new_n1109_ & new_n996_;
  assign new_n1262_ = ~new_n1183_ | ~new_n553_;
  assign new_n1263_ = ~new_n1110_;
  assign new_n1264_ = new_n1111_;
  assign new_n1265_ = ~new_n1184_ | ~new_n554_;
  assign new_n1266_ = new_n1112_;
  assign new_n1267_ = ~new_n1113_;
  assign new_n1268_ = new_n1114_ & new_n999_;
  assign new_n1269_ = new_n1115_ & new_n1001_;
  assign new_n1270_ = ~new_n1187_ | ~new_n557_;
  assign new_n1271_ = new_n1116_ & new_n1189_ & new_n1197_;
  assign new_n1272_ = new_n1189_ & new_n1116_;
  assign new_n1273_ = new_n1189_ & new_n1116_;
  assign new_n1274_ = ~new_n1188_ | ~new_n558_;
  assign new_n1275_ = new_n1191_ & new_n1117_;
  assign new_n1276_ = new_n1117_ & new_n1191_ & new_n1198_;
  assign new_n1277_ = new_n1191_ & new_n1117_;
  assign new_n1278_ = new_n1118_ & new_n1002_;
  assign new_n1279_ = new_n1119_ & new_n1004_;
  assign new_n1280_ = ~new_n1229_ | ~new_n561_;
  assign new_n1281_ = ~new_n1230_ | ~new_n562_;
  assign new_n1282_ = new_n1122_ & new_n1007_;
  assign new_n1283_ = new_n1123_ & new_n1009_;
  assign new_n1284_ = ~new_n1232_ | ~new_n565_;
  assign new_n1285_ = ~new_n1233_ | ~new_n566_;
  assign new_n1286_ = ~new_n1127_;
  assign new_n1287_ = ~new_n1129_;
  assign new_n1288_ = ~new_n1236_ | ~new_n567_;
  assign new_n1289_ = ~new_n1237_ | ~new_n568_;
  assign new_n1290_ = new_n1132_ & new_n1012_;
  assign new_n1291_ = new_n1133_ & new_n1014_;
  assign new_n1292_ = ~new_n1223_ | ~new_n571_;
  assign new_n1293_ = ~new_n1222_ | ~new_n572_;
  assign new_n1294_ = new_n1136_ & new_n1017_;
  assign new_n1295_ = new_n1137_ & new_n1019_;
  assign new_n1296_ = ~new_n1226_ | ~new_n575_;
  assign new_n1297_ = new_n1138_;
  assign new_n1298_ = ~new_n1139_;
  assign new_n1299_ = ~new_n1225_ | ~new_n576_;
  assign new_n1300_ = ~new_n1140_;
  assign new_n1301_ = new_n1141_;
  assign new_n1302_ = new_n1142_ & new_n1021_;
  assign new_n1303_ = new_n1143_ & new_n1023_;
  assign new_n1304_ = ~new_n1211_ | ~new_n579_;
  assign new_n1305_ = ~new_n1210_ | ~new_n580_;
  assign new_n1306_ = new_n1146_ & new_n1024_;
  assign new_n1307_ = new_n1147_ & new_n1026_;
  assign new_n1308_ = ~new_n1215_ | ~new_n583_;
  assign new_n1309_ = ~new_n1214_ | ~new_n584_;
  assign new_n1310_ = new_n1150_ & new_n1029_;
  assign new_n1311_ = new_n1151_ & new_n1031_;
  assign new_n1312_ = ~new_n1218_ | ~new_n587_;
  assign new_n1313_ = ~new_n1217_ | ~new_n588_;
  assign new_n1314_ = new_n1154_ & new_n1032_;
  assign new_n1315_ = new_n1155_ & new_n1034_;
  assign new_n1316_ = ~new_n1208_ | ~new_n592_;
  assign new_n1317_ = ~new_n1156_;
  assign new_n1318_ = new_n1157_;
  assign new_n1319_ = ~new_n1207_ | ~new_n593_;
  assign new_n1320_ = ~new_n1165_ | ~new_n1159_;
  assign new_n1321_ = new_n1161_;
  assign new_n1322_ = new_n1163_;
  assign new_n1323_ = new_n1164_;
  assign new_n1324_ = new_n1164_;
  assign new_n1325_ = ~new_n1165_;
  assign new_n1326_ = ~new_n1167_;
  assign new_n1327_ = ~new_n1167_;
  assign new_n1328_ = ~new_n1168_;
  assign new_n1329_ = ~new_n1169_;
  assign new_n1330_ = ~new_n1170_;
  assign new_n1331_ = ~new_n1172_;
  assign new_n1332_ = ~new_n1173_;
  assign new_n1333_ = ~new_n1174_;
  assign new_n1334_ = ~new_n1178_ | ~new_n1177_;
  assign new_n1335_ = ~new_n1178_;
  assign new_n1336_ = ~new_n1179_;
  assign new_n1337_ = ~new_n1180_;
  assign new_n1338_ = new_n627_ & new_n1171_ & new_n1160_;
  assign new_n1339_ = new_n849_ & new_n1037_ & new_n1171_;
  assign new_n1340_ = new_n850_ & new_n1160_ & new_n1042_;
  assign new_n1341_ = ~new_n1182_;
  assign new_n1342_ = ~new_n1183_;
  assign new_n1343_ = ~new_n1184_;
  assign new_n1344_ = ~new_n1049_ | ~new_n1195_;
  assign new_n1345_ = ~new_n1186_;
  assign new_n1346_ = ~new_n1187_;
  assign new_n1347_ = ~new_n1188_;
  assign new_n1348_ = new_n1189_;
  assign new_n1349_ = new_n1189_;
  assign new_n1350_ = new_n1197_ & new_n1190_;
  assign new_n1351_ = new_n1191_;
  assign new_n1352_ = new_n1191_;
  assign new_n1353_ = new_n1198_ & new_n1192_;
  assign new_n1354_ = ~new_n1193_;
  assign new_n1355_ = ~new_n1194_ | ~new_n1201_;
  assign new_n1356_ = ~new_n1194_;
  assign new_n1357_ = ~new_n1053_ | ~new_n1185_;
  assign new_n1358_ = ~new_n1196_;
  assign new_n1359_ = new_n1197_;
  assign new_n1360_ = new_n1197_;
  assign new_n1361_ = new_n1198_;
  assign new_n1362_ = new_n1198_;
  assign new_n1363_ = ~new_n1199_;
  assign new_n1364_ = ~new_n1200_;
  assign new_n1365_ = ~new_n1235_ | ~new_n1204_;
  assign new_n1366_ = new_n1219_ & new_n1062_ & new_n1059_;
  assign new_n1367_ = new_n1220_ & new_n1212_ & new_n1205_;
  assign new_n1368_ = ~new_n1206_;
  assign new_n1369_ = ~new_n1207_;
  assign new_n1370_ = ~new_n1208_;
  assign new_n1371_ = ~new_n1209_;
  assign new_n1372_ = ~new_n1210_;
  assign new_n1373_ = ~new_n1211_;
  assign new_n1374_ = ~new_n1213_;
  assign new_n1375_ = ~new_n1214_;
  assign new_n1376_ = ~new_n1215_;
  assign new_n1377_ = ~new_n1216_;
  assign new_n1378_ = ~new_n1217_;
  assign new_n1379_ = ~new_n1218_;
  assign new_n1380_ = ~new_n1219_;
  assign new_n1381_ = ~new_n1220_;
  assign new_n1382_ = ~new_n1221_;
  assign new_n1383_ = ~new_n1222_;
  assign new_n1384_ = ~new_n1223_;
  assign new_n1385_ = ~new_n1224_;
  assign new_n1386_ = ~new_n1225_;
  assign new_n1387_ = ~new_n1226_;
  assign new_n1388_ = ~new_n1234_ | ~new_n1227_;
  assign new_n1389_ = ~new_n1228_;
  assign new_n1390_ = ~new_n1229_;
  assign new_n1391_ = ~new_n1230_;
  assign new_n1392_ = ~new_n1231_;
  assign new_n1393_ = ~new_n1232_;
  assign new_n1394_ = ~new_n1233_;
  assign new_n1395_ = ~new_n1234_;
  assign new_n1396_ = ~new_n1235_;
  assign new_n1397_ = ~new_n1236_;
  assign new_n1398_ = ~new_n1237_;
  assign po039 = new_n1089_ & new_n744_;
  assign po040 = new_n1090_ & new_n744_;
  assign po041 = new_n1088_ & new_n744_;
  assign po042 = new_n1091_ & new_n744_;
  assign new_n1403_ = pi020 & new_n1161_;
  assign po035 = ~new_n1238_;
  assign po036 = ~new_n1239_;
  assign po037 = ~new_n1240_;
  assign po038 = ~new_n1241_;
  assign new_n1408_ = new_n490_ & new_n1256_ & new_n497_;
  assign new_n1409_ = new_n490_ & new_n1261_ & new_n497_;
  assign new_n1410_ = new_n490_ & new_n1268_ & new_n497_;
  assign new_n1411_ = new_n491_ & new_n1291_ & new_n498_;
  assign new_n1412_ = new_n491_ & new_n1295_ & new_n498_;
  assign new_n1413_ = new_n491_ & new_n1279_ & new_n498_;
  assign new_n1414_ = new_n491_ & new_n1283_ & new_n498_;
  assign new_n1415_ = new_n493_ & new_n1247_ & new_n499_;
  assign new_n1416_ = new_n493_ & new_n1250_ & new_n499_;
  assign new_n1417_ = new_n495_ & new_n1315_ & new_n500_;
  assign new_n1418_ = new_n495_ & new_n1302_ & new_n500_;
  assign new_n1419_ = new_n495_ & new_n1307_ & new_n500_;
  assign new_n1420_ = new_n495_ & new_n1310_ & new_n500_;
  assign new_n1421_ = ~new_n1246_;
  assign new_n1422_ = ~new_n1247_;
  assign new_n1423_ = ~new_n350_ | ~new_n1329_;
  assign new_n1424_ = ~new_n351_ | ~new_n1328_;
  assign new_n1425_ = ~new_n1250_;
  assign new_n1426_ = ~new_n1251_;
  assign new_n1427_ = ~new_n352_ | ~new_n1333_;
  assign new_n1428_ = ~new_n353_ | ~new_n1332_;
  assign new_n1429_ = ~new_n1257_ | ~new_n1100_;
  assign new_n1430_ = ~new_n1102_ | ~new_n1254_;
  assign new_n1431_ = ~new_n1255_ | ~new_n1103_;
  assign new_n1432_ = ~new_n1256_;
  assign new_n1433_ = ~new_n1257_;
  assign new_n1434_ = ~new_n356_ | ~new_n1337_;
  assign new_n1435_ = ~new_n357_ | ~new_n1336_;
  assign new_n1436_ = ~new_n1260_;
  assign new_n1437_ = ~new_n1261_;
  assign new_n1438_ = ~new_n358_ | ~new_n1342_;
  assign new_n1439_ = ~new_n1264_;
  assign new_n1440_ = ~new_n359_ | ~new_n1343_;
  assign new_n1441_ = ~new_n1266_;
  assign new_n1442_ = ~new_n1268_;
  assign new_n1443_ = ~new_n1269_;
  assign new_n1444_ = ~new_n360_ | ~new_n1346_;
  assign new_n1445_ = ~new_n361_ | ~new_n1347_;
  assign new_n1446_ = ~new_n1278_;
  assign new_n1447_ = ~new_n1279_;
  assign new_n1448_ = ~new_n362_ | ~new_n1390_;
  assign new_n1449_ = ~new_n363_ | ~new_n1391_;
  assign new_n1450_ = ~new_n1282_;
  assign new_n1451_ = ~new_n1283_;
  assign new_n1452_ = ~new_n364_ | ~new_n1393_;
  assign new_n1453_ = ~new_n365_ | ~new_n1394_;
  assign new_n1454_ = new_n1286_ & new_n1126_;
  assign new_n1455_ = new_n1287_ & new_n1128_;
  assign new_n1456_ = ~new_n366_ | ~new_n1397_;
  assign new_n1457_ = ~new_n367_ | ~new_n1398_;
  assign new_n1458_ = ~new_n1290_;
  assign new_n1459_ = ~new_n1291_;
  assign new_n1460_ = ~new_n368_ | ~new_n1384_;
  assign new_n1461_ = ~new_n369_ | ~new_n1383_;
  assign new_n1462_ = ~new_n1294_;
  assign new_n1463_ = ~new_n1295_;
  assign new_n1464_ = ~new_n370_ | ~new_n1387_;
  assign new_n1465_ = ~new_n1297_;
  assign new_n1466_ = ~new_n371_ | ~new_n1386_;
  assign new_n1467_ = ~new_n1301_;
  assign new_n1468_ = ~new_n1302_;
  assign new_n1469_ = ~new_n1303_;
  assign new_n1470_ = ~new_n372_ | ~new_n1373_;
  assign new_n1471_ = ~new_n373_ | ~new_n1372_;
  assign new_n1472_ = ~new_n1306_;
  assign new_n1473_ = ~new_n1307_;
  assign new_n1474_ = ~new_n374_ | ~new_n1376_;
  assign new_n1475_ = ~new_n375_ | ~new_n1375_;
  assign new_n1476_ = ~new_n1310_;
  assign new_n1477_ = ~new_n1311_;
  assign new_n1478_ = ~new_n376_ | ~new_n1379_;
  assign new_n1479_ = ~new_n377_ | ~new_n1378_;
  assign new_n1480_ = ~new_n1314_;
  assign new_n1481_ = ~new_n1315_;
  assign new_n1482_ = ~new_n380_ | ~new_n1370_;
  assign new_n1483_ = ~new_n1318_;
  assign new_n1484_ = ~new_n381_ | ~new_n1369_;
  assign new_n1485_ = ~new_n1036_ | ~new_n1325_;
  assign new_n1486_ = ~new_n1321_;
  assign new_n1487_ = new_n1162_ | new_n1403_;
  assign new_n1488_ = ~new_n1322_;
  assign new_n1489_ = ~new_n1323_;
  assign new_n1490_ = ~new_n1324_;
  assign new_n1491_ = ~new_n1327_;
  assign new_n1492_ = ~new_n1170_ | ~new_n1331_;
  assign new_n1493_ = ~new_n1172_ | ~new_n1330_;
  assign new_n1494_ = ~new_n1046_ | ~new_n1335_;
  assign new_n1495_ = ~new_n1339_ & ~new_n1338_;
  assign new_n1496_ = ~new_n1340_ & ~new_n1181_;
  assign new_n1497_ = ~new_n1182_ | ~new_n1345_;
  assign new_n1498_ = ~new_n1344_ | ~new_n1357_;
  assign new_n1499_ = ~new_n1186_ | ~new_n1341_;
  assign new_n1500_ = ~new_n1348_;
  assign new_n1501_ = ~new_n1349_;
  assign new_n1502_ = ~new_n1351_;
  assign new_n1503_ = ~new_n1352_;
  assign new_n1504_ = ~new_n1193_ | ~new_n1363_;
  assign new_n1505_ = ~new_n1359_;
  assign new_n1506_ = ~new_n1360_;
  assign new_n1507_ = ~new_n1361_;
  assign new_n1508_ = ~new_n1362_;
  assign new_n1509_ = ~new_n1199_ | ~new_n1354_;
  assign new_n1510_ = new_n1364_ & new_n1200_;
  assign new_n1511_ = ~new_n1056_ | ~new_n1356_;
  assign new_n1512_ = ~new_n1058_ | ~new_n1396_;
  assign new_n1513_ = new_n1381_ & new_n1059_ & new_n1212_;
  assign new_n1514_ = ~new_n1206_ | ~new_n1371_;
  assign new_n1515_ = ~new_n1209_ | ~new_n1368_;
  assign new_n1516_ = new_n1380_ & new_n1205_ & new_n1062_;
  assign new_n1517_ = ~new_n1213_ | ~new_n1377_;
  assign new_n1518_ = ~new_n1216_ | ~new_n1374_;
  assign new_n1519_ = ~new_n1221_ | ~new_n1385_;
  assign new_n1520_ = ~new_n1224_ | ~new_n1382_;
  assign new_n1521_ = ~new_n1070_ | ~new_n1395_;
  assign new_n1522_ = ~new_n1228_ | ~new_n1392_;
  assign new_n1523_ = ~new_n1231_ | ~new_n1389_;
  assign new_n1524_ = ~new_n1321_ | ~new_n772_;
  assign new_n1525_ = new_n491_ & new_n1454_ & new_n498_;
  assign new_n1526_ = ~new_n1246_ | ~new_n1426_;
  assign new_n1527_ = ~new_n1248_ | ~new_n1423_;
  assign new_n1528_ = ~new_n1424_ | ~new_n1249_;
  assign new_n1529_ = ~new_n1251_ | ~new_n1421_;
  assign new_n1530_ = ~new_n1427_ | ~new_n1252_;
  assign new_n1531_ = new_n1431_ & new_n1098_;
  assign new_n1532_ = ~new_n1253_ | ~new_n1428_;
  assign new_n1533_ = new_n1430_ & new_n1099_;
  assign new_n1534_ = new_n1430_ & new_n1099_;
  assign new_n1535_ = ~new_n986_ | ~new_n1433_;
  assign new_n1536_ = new_n1432_ & new_n1101_ & new_n1422_ & new_n1425_;
  assign new_n1537_ = new_n1430_;
  assign new_n1538_ = new_n1430_;
  assign new_n1539_ = new_n1431_;
  assign new_n1540_ = ~new_n1258_ | ~new_n1434_;
  assign new_n1541_ = ~new_n1435_ | ~new_n1259_;
  assign new_n1542_ = ~new_n1260_ | ~new_n1443_;
  assign new_n1543_ = ~new_n1262_ | ~new_n1438_;
  assign new_n1544_ = ~new_n1440_ | ~new_n1265_;
  assign new_n1545_ = ~new_n1269_ | ~new_n1436_;
  assign new_n1546_ = ~new_n1444_ | ~new_n1270_;
  assign new_n1547_ = ~new_n1274_ | ~new_n1445_;
  assign new_n1548_ = ~new_n1278_ | ~new_n1462_;
  assign new_n1549_ = new_n1451_ & new_n1447_ & new_n1459_ & new_n1463_;
  assign new_n1550_ = ~new_n1448_ | ~new_n1280_;
  assign new_n1551_ = ~new_n1281_ | ~new_n1449_;
  assign new_n1552_ = ~new_n1284_ | ~new_n1452_;
  assign new_n1553_ = ~new_n1453_ | ~new_n1285_;
  assign new_n1554_ = ~new_n1455_;
  assign new_n1555_ = new_n1455_;
  assign new_n1556_ = ~new_n1456_ | ~new_n1288_;
  assign new_n1557_ = ~new_n1289_ | ~new_n1457_;
  assign new_n1558_ = ~new_n1290_ | ~new_n1477_;
  assign new_n1559_ = ~new_n1292_ | ~new_n1460_;
  assign new_n1560_ = ~new_n1461_ | ~new_n1293_;
  assign new_n1561_ = ~new_n1294_ | ~new_n1446_;
  assign new_n1562_ = ~new_n1464_ | ~new_n1296_;
  assign new_n1563_ = ~new_n1299_ | ~new_n1466_;
  assign new_n1564_ = new_n1476_ & new_n1473_ & new_n1481_ & new_n1468_;
  assign new_n1565_ = ~new_n1303_ | ~new_n1472_;
  assign new_n1566_ = ~new_n1470_ | ~new_n1304_;
  assign new_n1567_ = ~new_n1305_ | ~new_n1471_;
  assign new_n1568_ = ~new_n1306_ | ~new_n1469_;
  assign new_n1569_ = ~new_n1308_ | ~new_n1474_;
  assign new_n1570_ = ~new_n1475_ | ~new_n1309_;
  assign new_n1571_ = ~new_n1311_ | ~new_n1458_;
  assign new_n1572_ = ~new_n1478_ | ~new_n1312_;
  assign new_n1573_ = ~new_n1313_ | ~new_n1479_;
  assign new_n1574_ = ~new_n1480_;
  assign new_n1575_ = ~new_n1316_ | ~new_n1482_;
  assign new_n1576_ = ~new_n1484_ | ~new_n1319_;
  assign new_n1577_ = ~new_n1320_ | ~new_n1485_;
  assign new_n1578_ = ~new_n1487_;
  assign new_n1579_ = ~new_n1493_ | ~new_n1492_;
  assign new_n1580_ = ~new_n1494_ | ~new_n1334_;
  assign new_n1581_ = ~new_n1495_ | ~new_n1496_;
  assign new_n1582_ = ~new_n1497_ | ~new_n1499_;
  assign new_n1583_ = ~new_n1498_;
  assign new_n1584_ = ~new_n1504_ | ~new_n1509_;
  assign new_n1585_ = ~new_n1355_ | ~new_n1511_;
  assign new_n1586_ = new_n1364_ | new_n1510_;
  assign new_n1587_ = new_n1202_ & new_n1358_ & new_n1437_ & new_n1442_;
  assign new_n1588_ = ~new_n1365_ | ~new_n1512_;
  assign new_n1589_ = ~new_n1516_ & ~new_n1366_;
  assign new_n1590_ = ~new_n1513_ & ~new_n1367_;
  assign new_n1591_ = ~new_n1514_ | ~new_n1515_;
  assign new_n1592_ = ~new_n1517_ | ~new_n1518_;
  assign new_n1593_ = ~new_n1519_ | ~new_n1520_;
  assign new_n1594_ = ~new_n1521_ | ~new_n1388_;
  assign new_n1595_ = ~new_n1522_ | ~new_n1523_;
  assign new_n1596_ = ~new_n484_ | ~new_n1486_;
  assign new_n1597_ = ~new_n1526_ | ~new_n1529_;
  assign new_n1598_ = new_n1527_;
  assign new_n1599_ = new_n1527_;
  assign new_n1600_ = new_n1430_ & new_n1532_ & new_n1094_;
  assign new_n1601_ = new_n1430_ & new_n1532_ & new_n1094_;
  assign new_n1602_ = new_n1430_ & new_n1094_ & new_n1532_ & new_n1540_;
  assign new_n1603_ = new_n1532_ & new_n1094_;
  assign new_n1604_ = new_n1532_ & new_n1094_;
  assign new_n1605_ = new_n1431_ & new_n1530_ & new_n1095_;
  assign new_n1606_ = new_n1431_ & new_n1095_ & new_n1530_ & new_n1541_;
  assign new_n1607_ = new_n1095_ & new_n1530_;
  assign new_n1608_ = new_n1528_;
  assign new_n1609_ = new_n1530_;
  assign new_n1610_ = new_n1098_ & new_n1431_ & new_n1541_;
  assign new_n1611_ = new_n1532_;
  assign new_n1612_ = new_n1532_;
  assign new_n1613_ = new_n1099_ & new_n1430_ & new_n1540_;
  assign new_n1614_ = ~new_n1535_ | ~new_n1429_;
  assign new_n1615_ = ~new_n1537_;
  assign new_n1616_ = ~new_n1538_;
  assign new_n1617_ = new_n1540_ & new_n988_;
  assign new_n1618_ = ~new_n1539_;
  assign new_n1619_ = new_n1541_ & new_n989_;
  assign new_n1620_ = new_n1540_;
  assign new_n1621_ = new_n1540_;
  assign new_n1622_ = new_n1541_;
  assign new_n1623_ = ~new_n1542_ | ~new_n1545_;
  assign new_n1624_ = new_n1543_;
  assign new_n1625_ = new_n1543_ & new_n1547_;
  assign new_n1626_ = new_n1543_;
  assign new_n1627_ = new_n1191_ & new_n1547_ & new_n1111_;
  assign new_n1628_ = new_n1191_ & new_n1111_ & new_n1547_ & new_n1198_;
  assign new_n1629_ = new_n1191_ & new_n1547_ & new_n1111_;
  assign new_n1630_ = new_n1547_ & new_n1111_;
  assign new_n1631_ = new_n1544_ & new_n1546_;
  assign new_n1632_ = ~new_n1544_;
  assign new_n1633_ = new_n1189_ & new_n1112_ & new_n1546_ & new_n1197_;
  assign new_n1634_ = new_n1189_ & new_n1112_ & new_n1546_;
  assign new_n1635_ = new_n1189_ & new_n1546_ & new_n1112_;
  assign new_n1636_ = new_n1546_ & new_n1112_;
  assign new_n1637_ = new_n1546_ & new_n1112_;
  assign new_n1638_ = new_n1546_;
  assign new_n1639_ = new_n1546_;
  assign new_n1640_ = new_n1547_;
  assign new_n1641_ = new_n1547_;
  assign new_n1642_ = ~new_n1561_ | ~new_n1548_;
  assign po044 = new_n1554_ & new_n1549_ & new_n1564_;
  assign new_n1644_ = new_n1550_;
  assign new_n1645_ = new_n1550_;
  assign new_n1646_ = new_n1556_ & new_n1550_ & new_n1553_ & new_n1562_;
  assign new_n1647_ = new_n1553_ & new_n1562_ & new_n1550_;
  assign new_n1648_ = new_n1562_ & new_n1550_;
  assign new_n1649_ = new_n1120_ & new_n1553_ & new_n1556_;
  assign new_n1650_ = new_n1553_ & new_n1120_;
  assign new_n1651_ = new_n1553_ & new_n1120_;
  assign new_n1652_ = new_n1563_ & new_n1551_;
  assign new_n1653_ = new_n1551_;
  assign new_n1654_ = new_n1557_ & new_n1552_ & new_n1563_ & new_n1551_;
  assign new_n1655_ = new_n1552_ & new_n1563_ & new_n1551_;
  assign new_n1656_ = new_n1551_;
  assign new_n1657_ = new_n1552_ & new_n1121_;
  assign new_n1658_ = new_n1121_ & new_n1552_ & new_n1557_;
  assign new_n1659_ = new_n1552_ & new_n1121_;
  assign new_n1660_ = ~new_n1555_ | ~new_n1450_;
  assign new_n1661_ = new_n1552_;
  assign new_n1662_ = new_n1552_;
  assign new_n1663_ = new_n1557_ & new_n1124_;
  assign new_n1664_ = new_n1553_;
  assign new_n1665_ = new_n1553_;
  assign new_n1666_ = new_n1556_ & new_n1125_;
  assign new_n1667_ = ~new_n1555_;
  assign new_n1668_ = new_n1556_;
  assign new_n1669_ = new_n1556_;
  assign new_n1670_ = new_n1557_;
  assign new_n1671_ = new_n1557_;
  assign new_n1672_ = ~new_n1571_ | ~new_n1558_;
  assign new_n1673_ = new_n1559_;
  assign new_n1674_ = new_n1559_;
  assign new_n1675_ = new_n1559_ & new_n1573_ & new_n1569_ & new_n1575_ & new_n1567_;
  assign new_n1676_ = new_n1566_ & new_n1560_ & new_n1570_ & new_n1572_ & new_n1576_;
  assign new_n1677_ = new_n1560_;
  assign new_n1678_ = ~new_n1562_;
  assign new_n1679_ = new_n1553_ & new_n1138_ & new_n1550_ & new_n1556_;
  assign new_n1680_ = new_n1553_ & new_n1138_ & new_n1550_;
  assign new_n1681_ = new_n1553_ & new_n1550_ & new_n1138_;
  assign new_n1682_ = new_n1550_ & new_n1138_;
  assign new_n1683_ = new_n1550_ & new_n1138_;
  assign new_n1684_ = new_n1563_;
  assign new_n1685_ = new_n1563_;
  assign new_n1686_ = new_n1552_ & new_n1551_ & new_n1141_;
  assign new_n1687_ = new_n1552_ & new_n1141_ & new_n1551_ & new_n1557_;
  assign new_n1688_ = new_n1552_ & new_n1551_ & new_n1141_;
  assign new_n1689_ = new_n1551_ & new_n1141_;
  assign new_n1690_ = ~new_n1565_ | ~new_n1568_;
  assign new_n1691_ = new_n1572_ & new_n1570_ & new_n1144_;
  assign new_n1692_ = new_n1572_ & new_n1144_ & new_n1570_ & new_n1560_;
  assign new_n1693_ = new_n1144_ & new_n1570_;
  assign new_n1694_ = new_n1566_;
  assign new_n1695_ = new_n1567_;
  assign new_n1696_ = new_n1567_ & new_n1573_ & new_n1575_ & new_n1569_;
  assign new_n1697_ = new_n1567_ & new_n1575_ & new_n1569_;
  assign new_n1698_ = new_n1567_;
  assign new_n1699_ = new_n1575_ & new_n1567_;
  assign new_n1700_ = new_n1573_ & new_n1569_ & new_n1145_;
  assign new_n1701_ = new_n1573_ & new_n1569_ & new_n1145_;
  assign new_n1702_ = new_n1573_ & new_n1145_ & new_n1569_ & new_n1559_;
  assign new_n1703_ = new_n1569_ & new_n1145_;
  assign new_n1704_ = new_n1569_ & new_n1145_;
  assign new_n1705_ = new_n1569_;
  assign new_n1706_ = new_n1569_;
  assign new_n1707_ = new_n1573_ & new_n1148_;
  assign new_n1708_ = new_n1573_ & new_n1148_;
  assign new_n1709_ = new_n1148_ & new_n1573_ & new_n1559_;
  assign new_n1710_ = new_n1570_;
  assign new_n1711_ = new_n1572_ & new_n1149_;
  assign new_n1712_ = new_n1149_ & new_n1572_ & new_n1560_;
  assign new_n1713_ = new_n1572_;
  assign new_n1714_ = new_n1560_ & new_n1152_;
  assign new_n1715_ = new_n1573_;
  assign new_n1716_ = new_n1573_;
  assign new_n1717_ = new_n1559_ & new_n1153_;
  assign new_n1718_ = new_n1575_;
  assign new_n1719_ = new_n1575_;
  assign new_n1720_ = new_n1573_ & new_n1157_ & new_n1567_ & new_n1569_;
  assign new_n1721_ = new_n1573_ & new_n1157_ & new_n1559_ & new_n1567_ & new_n1569_;
  assign new_n1722_ = new_n1573_ & new_n1157_ & new_n1567_ & new_n1569_;
  assign new_n1723_ = new_n1157_ & new_n1567_ & new_n1569_;
  assign new_n1724_ = new_n1567_ & new_n1157_;
  assign new_n1725_ = new_n1157_ & new_n1567_ & new_n1569_;
  assign new_n1726_ = new_n1576_;
  assign new_n1727_ = new_n1572_ & new_n1158_ & new_n1566_ & new_n1570_;
  assign new_n1728_ = new_n1572_ & new_n1158_ & new_n1560_ & new_n1566_ & new_n1570_;
  assign new_n1729_ = new_n1566_ & new_n1158_;
  assign new_n1730_ = new_n1158_ & new_n1566_ & new_n1570_;
  assign new_n1731_ = ~new_n1577_;
  assign new_n1732_ = new_n1528_ & new_n1541_ & new_n1530_ & new_n1431_ & new_n1161_;
  assign new_n1733_ = new_n1431_ & new_n1162_ & new_n1528_ & new_n1530_;
  assign new_n1734_ = new_n1431_ & new_n1162_ & new_n1541_ & new_n1528_ & new_n1530_;
  assign new_n1735_ = new_n1528_ & new_n1162_;
  assign new_n1736_ = new_n1162_ & new_n1528_ & new_n1530_;
  assign new_n1737_ = new_n1430_ & new_n1163_ & new_n1527_ & new_n1532_;
  assign new_n1738_ = new_n1430_ & new_n1163_ & new_n1540_ & new_n1527_ & new_n1532_;
  assign new_n1739_ = new_n1430_ & new_n1163_ & new_n1527_ & new_n1532_;
  assign new_n1740_ = new_n1163_ & new_n1527_ & new_n1532_;
  assign new_n1741_ = new_n1527_ & new_n1163_;
  assign new_n1742_ = new_n1163_ & new_n1527_ & new_n1532_;
  assign new_n1743_ = new_n1540_ & new_n1430_ & new_n1532_ & new_n1164_ & new_n1527_;
  assign new_n1744_ = new_n1527_ & new_n1430_ & new_n1164_ & new_n1532_;
  assign new_n1745_ = new_n1164_ & new_n1527_;
  assign new_n1746_ = new_n1527_ & new_n1164_ & new_n1532_;
  assign po043 = new_n1326_ & new_n1587_ & new_n1536_;
  assign new_n1748_ = ~new_n1579_;
  assign new_n1749_ = new_n1580_;
  assign new_n1750_ = new_n1580_;
  assign new_n1751_ = ~new_n1581_ | ~new_n1583_;
  assign new_n1752_ = ~new_n1581_;
  assign new_n1753_ = ~new_n1582_;
  assign new_n1754_ = new_n1197_ & new_n1546_ & new_n1189_ & new_n1544_;
  assign new_n1755_ = new_n1189_ & new_n1544_ & new_n1546_;
  assign new_n1756_ = new_n1198_ & new_n1191_ & new_n1543_ & new_n1547_;
  assign new_n1757_ = new_n1191_ & new_n1543_ & new_n1547_;
  assign new_n1758_ = ~new_n1584_;
  assign new_n1759_ = ~new_n1585_;
  assign new_n1760_ = new_n1588_;
  assign new_n1761_ = new_n1588_;
  assign new_n1762_ = ~new_n1590_ | ~new_n1589_;
  assign new_n1763_ = ~new_n1591_;
  assign new_n1764_ = ~new_n1592_;
  assign new_n1765_ = ~new_n1593_;
  assign new_n1766_ = ~new_n1594_;
  assign new_n1767_ = ~new_n1595_;
  assign new_n1768_ = ~new_n1586_ | ~pi060;
  assign new_n1769_ = new_n1431_ & new_n1528_ & new_n1530_ & pi020 & new_n1161_;
  assign new_n1770_ = new_n1528_ & pi020 & new_n1161_;
  assign new_n1771_ = ~new_n1524_ | ~new_n1596_;
  assign new_n1772_ = new_n1528_ & new_n1530_ & pi020 & new_n1161_;
  assign new_n1773_ = new_n1572_ & new_n1566_ & new_n1570_ & pi001 & new_n1576_;
  assign new_n1774_ = pi001 & new_n1576_;
  assign new_n1775_ = new_n1566_ & pi001 & new_n1576_;
  assign new_n1776_ = new_n1566_ & new_n1570_ & pi001 & new_n1576_;
  assign new_n1777_ = new_n493_ & new_n1771_ & new_n309_;
  assign new_n1778_ = ~new_n1597_;
  assign new_n1779_ = ~new_n1598_;
  assign new_n1780_ = ~new_n1599_;
  assign new_n1781_ = new_n1094_ | new_n1741_;
  assign new_n1782_ = new_n1770_ | new_n1095_ | new_n1735_;
  assign new_n1783_ = ~new_n1608_;
  assign new_n1784_ = ~new_n1609_;
  assign new_n1785_ = new_n1772_ | new_n1736_ | new_n1098_ | new_n1607_;
  assign new_n1786_ = ~new_n1611_;
  assign new_n1787_ = ~new_n1612_;
  assign new_n1788_ = ~new_n1742_ & ~new_n1099_ & ~new_n1603_;
  assign new_n1789_ = new_n1746_ | new_n1740_ | new_n1099_ | new_n1604_;
  assign new_n1790_ = new_n1614_;
  assign new_n1791_ = new_n1614_;
  assign new_n1792_ = ~new_n1739_ & ~new_n1600_ & ~new_n988_ & ~new_n1533_;
  assign new_n1793_ = new_n1744_ | new_n1737_ | new_n1601_ | new_n988_ | new_n1534_;
  assign new_n1794_ = new_n1769_ | new_n1733_ | new_n1605_ | new_n989_ | new_n1531_;
  assign new_n1795_ = ~new_n1620_;
  assign new_n1796_ = ~new_n1621_;
  assign new_n1797_ = new_n1738_ | new_n1602_ | new_n1613_ | new_n1106_ | new_n1617_;
  assign new_n1798_ = ~new_n1622_;
  assign new_n1799_ = new_n1734_ | new_n1606_ | new_n1610_ | new_n1107_ | new_n1619_;
  assign new_n1800_ = ~new_n1623_ | ~new_n1759_;
  assign new_n1801_ = ~new_n1623_;
  assign new_n1802_ = ~new_n1624_;
  assign new_n1803_ = ~new_n1626_;
  assign new_n1804_ = ~new_n1638_ | ~new_n1441_;
  assign new_n1805_ = ~new_n1639_ | ~new_n1267_;
  assign new_n1806_ = ~new_n1638_;
  assign new_n1807_ = ~new_n1639_;
  assign new_n1808_ = ~new_n1116_ & ~new_n1637_;
  assign new_n1809_ = new_n1631_ | new_n1116_ | new_n1636_;
  assign new_n1810_ = ~new_n1640_;
  assign new_n1811_ = ~new_n1641_;
  assign new_n1812_ = new_n1117_ | new_n1630_;
  assign new_n1813_ = ~new_n1642_;
  assign new_n1814_ = ~new_n1644_;
  assign new_n1815_ = ~new_n1645_;
  assign po048 = new_n1646_ & new_n1676_;
  assign new_n1817_ = ~new_n1120_ & ~new_n1683_;
  assign new_n1818_ = new_n1648_ | new_n1120_ | new_n1682_;
  assign new_n1819_ = ~new_n1653_;
  assign po045 = new_n1654_ & new_n1675_;
  assign new_n1821_ = ~new_n1656_;
  assign new_n1822_ = new_n1121_ | new_n1689_;
  assign new_n1823_ = ~new_n1282_ | ~new_n1667_;
  assign new_n1824_ = ~new_n1661_;
  assign new_n1825_ = ~new_n1662_;
  assign new_n1826_ = ~new_n1688_ & ~new_n1124_ & ~new_n1657_;
  assign new_n1827_ = new_n1655_ | new_n1686_ | new_n1124_ | new_n1659_;
  assign new_n1828_ = ~new_n1664_;
  assign new_n1829_ = ~new_n1665_;
  assign new_n1830_ = ~new_n1680_ & ~new_n1125_ & ~new_n1651_;
  assign new_n1831_ = new_n1647_ | new_n1681_ | new_n1125_ | new_n1650_;
  assign new_n1832_ = ~new_n1668_;
  assign new_n1833_ = ~new_n1669_;
  assign new_n1834_ = new_n1679_ | new_n1649_ | new_n1130_ | new_n1666_;
  assign new_n1835_ = new_n1687_ | new_n1658_ | new_n1131_ | new_n1663_;
  assign new_n1836_ = ~new_n1670_;
  assign new_n1837_ = ~new_n1671_;
  assign new_n1838_ = new_n1672_;
  assign new_n1839_ = new_n1672_;
  assign new_n1840_ = ~new_n1673_;
  assign new_n1841_ = ~new_n1674_;
  assign new_n1842_ = ~new_n1675_;
  assign new_n1843_ = new_n1721_ | new_n1702_ | new_n1709_ | new_n1134_ | new_n1717_;
  assign new_n1844_ = ~new_n1677_;
  assign new_n1845_ = new_n1728_ | new_n1692_ | new_n1712_ | new_n1135_ | new_n1714_;
  assign new_n1846_ = ~new_n1644_ | ~new_n1465_;
  assign new_n1847_ = ~new_n1645_ | ~new_n1298_;
  assign new_n1848_ = ~new_n1684_;
  assign new_n1849_ = ~new_n1685_;
  assign new_n1850_ = ~new_n1690_;
  assign new_n1851_ = new_n1775_ | new_n1144_ | new_n1729_;
  assign new_n1852_ = ~new_n1694_;
  assign new_n1853_ = ~new_n1695_;
  assign new_n1854_ = ~new_n1698_;
  assign new_n1855_ = new_n1145_ | new_n1724_;
  assign new_n1856_ = ~new_n1705_;
  assign new_n1857_ = ~new_n1706_;
  assign new_n1858_ = ~new_n1725_ & ~new_n1148_ & ~new_n1703_;
  assign new_n1859_ = new_n1697_ | new_n1723_ | new_n1148_ | new_n1704_;
  assign new_n1860_ = ~new_n1710_;
  assign new_n1861_ = new_n1776_ | new_n1730_ | new_n1149_ | new_n1693_;
  assign new_n1862_ = ~new_n1713_;
  assign new_n1863_ = new_n1773_ | new_n1727_ | new_n1691_ | new_n1152_ | new_n1711_;
  assign new_n1864_ = ~new_n1715_;
  assign new_n1865_ = ~new_n1716_;
  assign new_n1866_ = ~new_n1722_ & ~new_n1700_ & ~new_n1153_ & ~new_n1707_;
  assign new_n1867_ = new_n1696_ | new_n1720_ | new_n1701_ | new_n1153_ | new_n1708_;
  assign new_n1868_ = ~new_n1718_;
  assign new_n1869_ = ~new_n1719_;
  assign new_n1870_ = ~new_n1726_;
  assign new_n1871_ = new_n1158_ | new_n1774_;
  assign new_n1872_ = new_n1750_ & new_n1577_ & new_n1579_;
  assign new_n1873_ = new_n1749_ & new_n1731_ & new_n1748_;
  assign po046 = new_n1754_ & new_n1732_;
  assign new_n1875_ = ~new_n1608_ | ~new_n1578_;
  assign po047 = new_n1756_ & new_n1743_;
  assign new_n1877_ = ~new_n1743_;
  assign new_n1878_ = ~new_n1749_;
  assign new_n1879_ = ~new_n1750_;
  assign new_n1880_ = ~new_n1582_ | ~new_n1758_;
  assign new_n1881_ = ~new_n1498_ | ~new_n1752_;
  assign new_n1882_ = ~new_n1634_ & ~new_n1190_ & ~new_n1273_;
  assign new_n1883_ = new_n1755_ | new_n1635_ | new_n1190_ | new_n1272_;
  assign new_n1884_ = ~new_n1629_ & ~new_n1192_ & ~new_n1275_;
  assign new_n1885_ = new_n1757_ | new_n1627_ | new_n1192_ | new_n1277_;
  assign new_n1886_ = ~new_n1584_ | ~new_n1753_;
  assign new_n1887_ = new_n1633_ | new_n1271_ | new_n1055_ | new_n1350_;
  assign new_n1888_ = new_n1628_ | new_n1276_ | new_n1055_ | new_n1353_;
  assign new_n1889_ = new_n1586_ & new_n1768_;
  assign new_n1890_ = ~new_n1760_;
  assign new_n1891_ = new_n1761_ & new_n1767_ & new_n1765_;
  assign new_n1892_ = ~new_n1761_;
  assign new_n1893_ = ~new_n1762_ | ~new_n1766_;
  assign new_n1894_ = ~new_n1762_;
  assign new_n1895_ = ~new_n1591_ | ~new_n1764_;
  assign new_n1896_ = ~new_n1592_ | ~new_n1763_;
  assign new_n1897_ = new_n1760_ & new_n1595_ & new_n1593_;
  assign new_n1898_ = new_n1768_ & pi060;
  assign new_n1899_ = new_n1732_ & pi020;
  assign new_n1900_ = ~new_n1771_;
  assign new_n1901_ = new_n1676_ & pi001;
  assign new_n1902_ = ~new_n1726_ | ~new_n786_;
  assign new_n1903_ = ~new_n1781_;
  assign new_n1904_ = ~new_n1782_ | ~new_n1784_;
  assign new_n1905_ = ~new_n1782_;
  assign new_n1906_ = ~new_n1785_;
  assign new_n1907_ = ~new_n1788_;
  assign new_n1908_ = ~new_n1789_;
  assign new_n1909_ = ~new_n1790_;
  assign new_n1910_ = ~new_n1791_;
  assign new_n1911_ = ~new_n1792_;
  assign new_n1912_ = ~new_n1793_;
  assign new_n1913_ = ~new_n1785_ | ~new_n1618_;
  assign new_n1914_ = ~new_n1794_ | ~new_n1798_;
  assign new_n1915_ = ~new_n1794_;
  assign new_n1916_ = ~new_n1797_;
  assign new_n1917_ = new_n1799_ | new_n1899_;
  assign new_n1918_ = new_n1812_ | new_n1625_;
  assign new_n1919_ = ~new_n1266_ | ~new_n1806_;
  assign new_n1920_ = ~new_n1113_ | ~new_n1807_;
  assign new_n1921_ = ~new_n1808_;
  assign new_n1922_ = ~new_n1809_;
  assign new_n1923_ = ~new_n1812_;
  assign new_n1924_ = new_n1845_ & new_n1646_;
  assign new_n1925_ = ~new_n1817_ | ~new_n1828_;
  assign new_n1926_ = ~new_n1817_;
  assign new_n1927_ = ~new_n1818_ | ~new_n1829_;
  assign new_n1928_ = ~new_n1818_;
  assign new_n1929_ = new_n1822_ | new_n1652_;
  assign new_n1930_ = new_n1654_ & new_n1843_;
  assign new_n1931_ = ~new_n1822_;
  assign new_n1932_ = ~new_n1823_ | ~new_n1660_;
  assign new_n1933_ = ~new_n1826_;
  assign new_n1934_ = ~new_n1827_;
  assign new_n1935_ = ~new_n1830_ | ~new_n1833_;
  assign new_n1936_ = ~new_n1830_;
  assign new_n1937_ = ~new_n1831_ | ~new_n1832_;
  assign new_n1938_ = ~new_n1831_;
  assign new_n1939_ = ~new_n1838_;
  assign new_n1940_ = ~new_n1839_;
  assign new_n1941_ = ~new_n1843_;
  assign new_n1942_ = ~new_n1863_ | ~new_n1844_;
  assign new_n1943_ = new_n1845_ | new_n1901_;
  assign new_n1944_ = ~new_n1297_ | ~new_n1814_;
  assign new_n1945_ = ~new_n1139_ | ~new_n1815_;
  assign new_n1946_ = ~new_n1851_ | ~new_n1860_;
  assign new_n1947_ = ~new_n1851_;
  assign new_n1948_ = ~new_n1871_ | ~new_n1852_;
  assign new_n1949_ = new_n1855_ | new_n1699_;
  assign new_n1950_ = ~new_n1855_;
  assign new_n1951_ = ~new_n1858_;
  assign new_n1952_ = ~new_n1859_;
  assign new_n1953_ = ~new_n1861_ | ~new_n1862_;
  assign new_n1954_ = ~new_n1861_;
  assign new_n1955_ = ~new_n1863_;
  assign new_n1956_ = ~new_n1866_;
  assign new_n1957_ = ~new_n1867_;
  assign new_n1958_ = new_n1839_ & new_n1690_ & new_n1480_;
  assign new_n1959_ = new_n1838_ & new_n1850_ & new_n1574_;
  assign new_n1960_ = ~new_n1859_ | ~new_n1317_;
  assign new_n1961_ = ~new_n1858_ | ~new_n1483_;
  assign new_n1962_ = ~new_n1871_;
  assign new_n1963_ = new_n1879_ & new_n1748_ & new_n1577_;
  assign new_n1964_ = ~new_n1487_ | ~new_n1783_;
  assign new_n1965_ = ~new_n1788_ | ~new_n1488_;
  assign new_n1966_ = new_n1781_ | new_n1745_;
  assign new_n1967_ = new_n1791_ & new_n1597_ & new_n1327_;
  assign new_n1968_ = new_n1790_ & new_n1778_ & new_n1491_;
  assign new_n1969_ = new_n1878_ & new_n1579_ & new_n1731_;
  assign new_n1970_ = ~new_n1881_ | ~new_n1751_;
  assign new_n1971_ = ~new_n1880_ | ~new_n1886_;
  assign new_n1972_ = ~new_n1808_ | ~new_n1500_;
  assign new_n1973_ = new_n1799_ & new_n1754_;
  assign new_n1974_ = ~new_n1809_ | ~new_n1501_;
  assign new_n1975_ = ~new_n1882_;
  assign new_n1976_ = ~new_n1883_;
  assign new_n1977_ = new_n1756_ & new_n1797_;
  assign new_n1978_ = ~new_n1884_;
  assign new_n1979_ = ~new_n1885_;
  assign new_n1980_ = ~new_n1585_ | ~new_n1801_;
  assign new_n1981_ = ~new_n1883_ | ~new_n1505_;
  assign new_n1982_ = ~new_n1882_ | ~new_n1506_;
  assign new_n1983_ = new_n1889_ | new_n1898_;
  assign new_n1984_ = ~new_n1895_ | ~new_n1896_;
  assign new_n1985_ = new_n1892_ & new_n1593_ & new_n1767_;
  assign new_n1986_ = ~new_n1594_ | ~new_n1894_;
  assign new_n1987_ = new_n1890_ & new_n1765_ & new_n1595_;
  assign new_n1988_ = new_n928_ | new_n1244_ | new_n1777_;
  assign new_n1989_ = ~new_n487_ | ~new_n1870_;
  assign new_n1990_ = new_n503_ & new_n1988_ & new_n505_;
  assign new_n1991_ = new_n509_ & new_n1988_ & new_n507_;
  assign new_n1992_ = new_n321_ & new_n1983_ & pi170;
  assign new_n1993_ = new_n523_ & new_n1988_ & new_n525_;
  assign new_n1994_ = new_n527_ & new_n1988_ & new_n529_;
  assign new_n1995_ = ~new_n1903_;
  assign new_n1996_ = ~new_n1609_ | ~new_n1905_;
  assign new_n1997_ = ~new_n1966_ | ~new_n1908_;
  assign new_n1998_ = ~new_n1539_ | ~new_n1906_;
  assign new_n1999_ = ~new_n1622_ | ~new_n1915_;
  assign new_n2000_ = ~new_n1917_;
  assign new_n2001_ = ~new_n1800_ | ~new_n1980_;
  assign new_n2002_ = ~new_n1918_;
  assign new_n2003_ = ~new_n1918_ | ~new_n1263_;
  assign new_n2004_ = ~new_n1923_ | ~new_n1439_;
  assign new_n2005_ = new_n1917_ & new_n1632_;
  assign new_n2006_ = ~new_n1804_ | ~new_n1919_;
  assign new_n2007_ = ~new_n1805_ | ~new_n1920_;
  assign new_n2008_ = ~new_n1923_;
  assign new_n2009_ = ~new_n1932_ | ~new_n1813_;
  assign new_n2010_ = ~new_n1929_;
  assign new_n2011_ = ~new_n1931_;
  assign new_n2012_ = ~new_n1932_;
  assign new_n2013_ = ~new_n1664_ | ~new_n1926_;
  assign new_n2014_ = ~new_n1665_ | ~new_n1928_;
  assign new_n2015_ = ~new_n1668_ | ~new_n1938_;
  assign new_n2016_ = ~new_n1669_ | ~new_n1936_;
  assign po053 = new_n1834_ | new_n1924_;
  assign po051 = new_n1835_ | new_n1930_;
  assign new_n2019_ = new_n1941_ & new_n1842_;
  assign new_n2020_ = ~new_n1677_ | ~new_n1955_;
  assign new_n2021_ = ~new_n1943_;
  assign new_n2022_ = new_n1943_ & new_n1678_;
  assign new_n2023_ = ~new_n1846_ | ~new_n1944_;
  assign new_n2024_ = ~new_n1847_ | ~new_n1945_;
  assign new_n2025_ = ~new_n1929_ | ~new_n1300_;
  assign new_n2026_ = ~new_n1931_ | ~new_n1467_;
  assign new_n2027_ = ~new_n1694_ | ~new_n1962_;
  assign new_n2028_ = ~new_n1949_;
  assign new_n2029_ = ~new_n1950_;
  assign new_n2030_ = ~new_n1710_ | ~new_n1947_;
  assign new_n2031_ = ~new_n1713_ | ~new_n1954_;
  assign new_n2032_ = new_n1939_ & new_n1480_ & new_n1850_;
  assign new_n2033_ = new_n1940_ & new_n1574_ & new_n1690_;
  assign new_n2034_ = ~new_n1156_ | ~new_n1952_;
  assign new_n2035_ = ~new_n1318_ | ~new_n1951_;
  assign new_n2036_ = ~new_n1963_ & ~new_n1872_;
  assign new_n2037_ = ~new_n1969_ & ~new_n1873_;
  assign new_n2038_ = ~new_n1875_ | ~new_n1964_;
  assign new_n2039_ = ~new_n1322_ | ~new_n1907_;
  assign new_n2040_ = new_n1916_ & new_n1877_;
  assign new_n2041_ = ~new_n1966_;
  assign new_n2042_ = new_n1909_ & new_n1327_ & new_n1778_;
  assign new_n2043_ = new_n1910_ & new_n1491_ & new_n1597_;
  assign po049 = new_n1970_;
  assign new_n2045_ = ~new_n1970_;
  assign new_n2046_ = ~new_n1971_;
  assign new_n2047_ = ~new_n1348_ | ~new_n1921_;
  assign new_n2048_ = ~new_n1349_ | ~new_n1922_;
  assign po052 = new_n1887_ | new_n1973_;
  assign po054 = new_n1888_ | new_n1977_;
  assign new_n2051_ = ~new_n1359_ | ~new_n1976_;
  assign new_n2052_ = ~new_n1360_ | ~new_n1975_;
  assign new_n2053_ = ~new_n1985_ & ~new_n1891_;
  assign new_n2054_ = ~new_n1986_ | ~new_n1893_;
  assign new_n2055_ = ~new_n1984_;
  assign new_n2056_ = ~new_n1987_ & ~new_n1897_;
  assign po055 = ~new_n1988_;
  assign new_n2058_ = ~new_n1902_ | ~new_n1989_;
  assign new_n2059_ = new_n493_ & new_n2038_ & new_n309_;
  assign new_n2060_ = new_n495_ & new_n2058_ & new_n310_;
  assign new_n2061_ = ~new_n1996_ | ~new_n1904_;
  assign new_n2062_ = ~new_n1789_ | ~new_n2041_;
  assign new_n2063_ = ~new_n1998_ | ~new_n1913_;
  assign new_n2064_ = ~new_n1999_ | ~new_n1914_;
  assign new_n2065_ = new_n2006_ & new_n2000_;
  assign new_n2066_ = ~new_n2001_;
  assign new_n2067_ = ~new_n1110_ | ~new_n2002_;
  assign new_n2068_ = ~new_n1264_ | ~new_n2008_;
  assign new_n2069_ = new_n1544_ & new_n2000_;
  assign new_n2070_ = ~new_n2007_;
  assign new_n2071_ = ~new_n1642_ | ~new_n2012_;
  assign new_n2072_ = ~new_n2013_ | ~new_n1925_;
  assign new_n2073_ = ~new_n2014_ | ~new_n1927_;
  assign new_n2074_ = ~new_n2016_ | ~new_n1935_;
  assign new_n2075_ = ~new_n2015_ | ~new_n1937_;
  assign new_n2076_ = ~new_n2019_;
  assign new_n2077_ = ~new_n2020_ | ~new_n1942_;
  assign new_n2078_ = new_n2023_ & new_n2021_;
  assign new_n2079_ = new_n1562_ & new_n2021_;
  assign new_n2080_ = ~new_n2024_;
  assign new_n2081_ = ~new_n1140_ | ~new_n2010_;
  assign new_n2082_ = ~new_n1301_ | ~new_n2011_;
  assign new_n2083_ = ~new_n2030_ | ~new_n1946_;
  assign new_n2084_ = ~new_n2027_ | ~new_n1948_;
  assign new_n2085_ = ~new_n2031_ | ~new_n1953_;
  assign new_n2086_ = ~new_n2033_ & ~new_n1958_;
  assign new_n2087_ = ~new_n2032_ & ~new_n1959_;
  assign new_n2088_ = ~new_n1960_ | ~new_n2034_;
  assign new_n2089_ = ~new_n1961_ | ~new_n2035_;
  assign new_n2090_ = ~new_n2037_ | ~new_n2036_;
  assign new_n2091_ = ~new_n2038_;
  assign new_n2092_ = ~new_n1965_ | ~new_n2039_;
  assign new_n2093_ = ~new_n2040_;
  assign new_n2094_ = ~new_n2043_ & ~new_n1967_;
  assign new_n2095_ = ~new_n2042_ & ~new_n1968_;
  assign new_n2096_ = ~new_n2047_ | ~new_n1972_;
  assign new_n2097_ = ~new_n2048_ | ~new_n1974_;
  assign new_n2098_ = ~new_n2051_ | ~new_n1981_;
  assign new_n2099_ = ~new_n2052_ | ~new_n1982_;
  assign new_n2100_ = ~new_n2053_ | ~new_n2056_;
  assign po050 = new_n2054_;
  assign new_n2102_ = ~new_n2054_;
  assign new_n2103_ = ~new_n2058_;
  assign new_n2104_ = new_n490_ & new_n2064_ & new_n307_;
  assign new_n2105_ = new_n491_ & new_n2077_ & new_n308_;
  assign new_n2106_ = new_n493_ & new_n2063_ & new_n309_;
  assign new_n2107_ = new_n493_ & new_n2061_ & new_n309_;
  assign new_n2108_ = new_n495_ & new_n2085_ & new_n310_;
  assign new_n2109_ = new_n495_ & new_n2083_ & new_n310_;
  assign new_n2110_ = new_n495_ & new_n2084_ & new_n310_;
  assign new_n2111_ = ~new_n2092_ | ~new_n1995_;
  assign new_n2112_ = ~new_n2061_;
  assign new_n2113_ = ~new_n1997_ | ~new_n2062_;
  assign new_n2114_ = ~new_n2063_;
  assign new_n2115_ = ~new_n2064_;
  assign new_n2116_ = new_n1917_ & new_n2097_;
  assign new_n2117_ = new_n1917_ & new_n2070_;
  assign new_n2118_ = new_n1917_ & new_n2098_;
  assign new_n2119_ = ~new_n2003_ | ~new_n2067_;
  assign new_n2120_ = ~new_n2004_ | ~new_n2068_;
  assign new_n2121_ = new_n2069_ | new_n2005_;
  assign new_n2122_ = ~new_n2071_ | ~new_n2009_;
  assign new_n2123_ = ~new_n2072_;
  assign new_n2124_ = ~new_n2074_;
  assign new_n2125_ = ~new_n2077_;
  assign new_n2126_ = new_n1943_ & new_n2073_;
  assign new_n2127_ = new_n1943_ & new_n2080_;
  assign new_n2128_ = new_n1943_ & new_n2075_;
  assign new_n2129_ = new_n2079_ | new_n2022_;
  assign new_n2130_ = ~new_n2025_ | ~new_n2081_;
  assign new_n2131_ = ~new_n2026_ | ~new_n2082_;
  assign new_n2132_ = ~new_n2083_;
  assign new_n2133_ = ~new_n2084_;
  assign new_n2134_ = ~new_n2088_ | ~new_n2028_;
  assign new_n2135_ = ~new_n2089_ | ~new_n2029_;
  assign new_n2136_ = ~new_n2085_;
  assign new_n2137_ = ~new_n2087_ | ~new_n2086_;
  assign new_n2138_ = ~new_n2088_;
  assign new_n2139_ = ~new_n2089_;
  assign new_n2140_ = ~new_n2090_;
  assign new_n2141_ = ~new_n2092_;
  assign new_n2142_ = ~new_n2095_ | ~new_n2094_;
  assign new_n2143_ = ~new_n2090_ | ~new_n2046_;
  assign new_n2144_ = ~new_n2096_;
  assign new_n2145_ = ~new_n2099_;
  assign new_n2146_ = ~new_n2100_;
  assign new_n2147_ = ~new_n2100_ | ~new_n2055_;
  assign new_n2148_ = new_n930_ | new_n1415_ | new_n2059_;
  assign new_n2149_ = new_n940_ | new_n1417_ | new_n2060_;
  assign new_n2150_ = new_n490_ & new_n2121_ & new_n307_;
  assign new_n2151_ = new_n491_ & new_n2129_ & new_n308_;
  assign new_n2152_ = new_n503_ & new_n2148_ & new_n505_;
  assign new_n2153_ = new_n503_ & new_n2149_ & new_n315_;
  assign new_n2154_ = new_n509_ & new_n2149_ & new_n317_;
  assign new_n2155_ = new_n509_ & new_n2148_ & new_n507_;
  assign new_n2156_ = new_n523_ & new_n2148_ & new_n525_;
  assign new_n2157_ = new_n523_ & new_n2149_ & new_n334_;
  assign new_n2158_ = new_n527_ & new_n2148_ & new_n529_;
  assign new_n2159_ = new_n527_ & new_n2149_ & new_n338_;
  assign new_n2160_ = ~new_n1903_ | ~new_n2141_;
  assign new_n2161_ = ~new_n2113_;
  assign new_n2162_ = ~new_n2113_ | ~new_n1912_;
  assign new_n2163_ = new_n2145_ & new_n2000_;
  assign new_n2164_ = new_n2065_ | new_n2117_;
  assign new_n2165_ = new_n2144_ & new_n2000_;
  assign new_n2166_ = ~new_n2142_ | ~new_n2066_;
  assign new_n2167_ = ~new_n2119_;
  assign new_n2168_ = ~new_n2120_;
  assign new_n2169_ = ~new_n2121_;
  assign new_n2170_ = ~new_n2122_;
  assign new_n2171_ = ~new_n2131_ | ~new_n1933_;
  assign new_n2172_ = ~new_n2130_ | ~new_n1934_;
  assign new_n2173_ = new_n2124_ & new_n2021_;
  assign new_n2174_ = new_n2078_ | new_n2127_;
  assign new_n2175_ = new_n2123_ & new_n2021_;
  assign new_n2176_ = ~new_n2129_;
  assign new_n2177_ = ~new_n2130_;
  assign new_n2178_ = ~new_n2131_;
  assign new_n2179_ = ~new_n1949_ | ~new_n2138_;
  assign new_n2180_ = ~new_n1950_ | ~new_n2139_;
  assign new_n2181_ = ~new_n2137_;
  assign new_n2182_ = ~new_n2142_;
  assign new_n2183_ = ~new_n1971_ | ~new_n2140_;
  assign new_n2184_ = ~new_n2120_ | ~new_n1978_;
  assign new_n2185_ = ~new_n2119_ | ~new_n1979_;
  assign new_n2186_ = ~new_n1984_ | ~new_n2146_;
  assign new_n2187_ = new_n929_ | new_n1087_ | new_n2106_;
  assign po056 = ~new_n2148_;
  assign new_n2189_ = new_n931_ | new_n1420_ | new_n2108_;
  assign new_n2190_ = new_n932_ | new_n1419_ | new_n2109_;
  assign new_n2191_ = new_n933_ | new_n1418_ | new_n2110_;
  assign new_n2192_ = new_n935_ | new_n1411_ | new_n2105_;
  assign new_n2193_ = new_n938_ | new_n1416_ | new_n2107_;
  assign po057 = ~new_n2149_;
  assign new_n2195_ = new_n961_ | new_n1408_ | new_n2104_;
  assign new_n2196_ = new_n490_ & new_n2164_ & new_n307_;
  assign new_n2197_ = new_n491_ & new_n2174_ & new_n308_;
  assign new_n2198_ = new_n502_ & new_n2195_ & new_n504_;
  assign new_n2199_ = new_n503_ & new_n2187_ & new_n505_;
  assign new_n2200_ = new_n503_ & new_n2193_ & new_n505_;
  assign new_n2201_ = new_n502_ & new_n2192_ & new_n314_;
  assign new_n2202_ = new_n503_ & new_n2189_ & new_n315_;
  assign new_n2203_ = new_n503_ & new_n2190_ & new_n315_;
  assign new_n2204_ = new_n503_ & new_n2191_ & new_n315_;
  assign new_n2205_ = new_n508_ & new_n2192_ & new_n316_;
  assign new_n2206_ = new_n508_ & new_n2195_ & new_n506_;
  assign new_n2207_ = new_n509_ & new_n2189_ & new_n317_;
  assign new_n2208_ = new_n509_ & new_n2190_ & new_n317_;
  assign new_n2209_ = new_n509_ & new_n2191_ & new_n317_;
  assign new_n2210_ = new_n509_ & new_n2187_ & new_n507_;
  assign new_n2211_ = new_n509_ & new_n2193_ & new_n507_;
  assign new_n2212_ = new_n523_ & new_n2193_ & new_n525_;
  assign new_n2213_ = new_n523_ & new_n2187_ & new_n525_;
  assign new_n2214_ = new_n524_ & new_n2195_ & new_n526_;
  assign new_n2215_ = new_n523_ & new_n2189_ & new_n334_;
  assign new_n2216_ = new_n523_ & new_n2190_ & new_n334_;
  assign new_n2217_ = new_n523_ & new_n2191_ & new_n334_;
  assign new_n2218_ = new_n524_ & new_n2192_ & new_n335_;
  assign new_n2219_ = new_n527_ & new_n2193_ & new_n529_;
  assign new_n2220_ = new_n527_ & new_n2187_ & new_n529_;
  assign new_n2221_ = new_n528_ & new_n2195_ & new_n530_;
  assign new_n2222_ = new_n527_ & new_n2189_ & new_n338_;
  assign new_n2223_ = new_n527_ & new_n2190_ & new_n338_;
  assign new_n2224_ = new_n527_ & new_n2191_ & new_n338_;
  assign new_n2225_ = new_n528_ & new_n2192_ & new_n339_;
  assign new_n2226_ = ~new_n2160_ | ~new_n2111_;
  assign new_n2227_ = ~new_n1793_ | ~new_n2161_;
  assign new_n2228_ = new_n2165_ | new_n2116_;
  assign new_n2229_ = new_n2163_ | new_n2118_;
  assign new_n2230_ = ~new_n2164_;
  assign new_n2231_ = ~new_n2001_ | ~new_n2182_;
  assign new_n2232_ = ~new_n2122_ | ~new_n2181_;
  assign new_n2233_ = ~new_n1826_ | ~new_n2178_;
  assign new_n2234_ = ~new_n1827_ | ~new_n2177_;
  assign new_n2235_ = new_n2175_ | new_n2126_;
  assign new_n2236_ = new_n2173_ | new_n2128_;
  assign new_n2237_ = ~new_n2174_;
  assign new_n2238_ = ~new_n2179_ | ~new_n2134_;
  assign new_n2239_ = ~new_n2180_ | ~new_n2135_;
  assign new_n2240_ = ~new_n2137_ | ~new_n2170_;
  assign new_n2241_ = ~new_n2183_ | ~new_n2143_;
  assign new_n2242_ = ~new_n1884_ | ~new_n2168_;
  assign new_n2243_ = ~new_n1885_ | ~new_n2167_;
  assign new_n2244_ = ~new_n2186_ | ~new_n2147_;
  assign new_n2245_ = new_n723_ | new_n921_ | new_n1994_ | new_n2159_;
  assign new_n2246_ = new_n724_ | new_n920_ | new_n1993_ | new_n2157_;
  assign po061 = ~new_n2187_;
  assign po065 = ~new_n2189_;
  assign po066 = ~new_n2190_;
  assign po067 = ~new_n2191_;
  assign po064 = ~new_n2192_;
  assign po062 = ~new_n2193_;
  assign new_n2253_ = new_n944_ | new_n1412_ | new_n2151_;
  assign new_n2254_ = new_n945_ | new_n1409_ | new_n2150_;
  assign po059 = new_n770_ | new_n972_ | new_n1991_ | new_n2154_;
  assign po063 = new_n771_ | new_n973_ | new_n1990_ | new_n2153_;
  assign po060 = ~new_n2195_;
  assign new_n2258_ = new_n490_ & new_n2229_ & new_n307_;
  assign new_n2259_ = new_n490_ & new_n2228_ & new_n307_;
  assign new_n2260_ = new_n491_ & new_n2236_ & new_n308_;
  assign new_n2261_ = new_n491_ & new_n2235_ & new_n308_;
  assign new_n2262_ = new_n502_ & new_n2254_ & new_n504_;
  assign new_n2263_ = new_n502_ & new_n2253_ & new_n314_;
  assign new_n2264_ = new_n508_ & new_n2253_ & new_n316_;
  assign new_n2265_ = new_n508_ & new_n2254_ & new_n506_;
  assign new_n2266_ = pi169 & new_n2229_ & pi170;
  assign new_n2267_ = new_n524_ & new_n2254_ & new_n526_;
  assign new_n2268_ = new_n524_ & new_n2253_ & new_n335_;
  assign new_n2269_ = new_n528_ & new_n2254_ & new_n530_;
  assign new_n2270_ = new_n528_ & new_n2253_ & new_n339_;
  assign new_n2271_ = ~new_n2226_;
  assign new_n2272_ = ~new_n2226_ | ~new_n1911_;
  assign new_n2273_ = ~new_n2227_ | ~new_n2162_;
  assign new_n2274_ = ~new_n2228_;
  assign new_n2275_ = ~new_n2229_;
  assign po058 = ~new_n2229_;
  assign new_n2277_ = ~new_n2231_ | ~new_n2166_;
  assign new_n2278_ = ~new_n2232_ | ~new_n2240_;
  assign new_n2279_ = ~new_n2233_ | ~new_n2171_;
  assign new_n2280_ = ~new_n2234_ | ~new_n2172_;
  assign new_n2281_ = ~new_n2235_;
  assign new_n2282_ = ~new_n2236_;
  assign new_n2283_ = ~new_n2238_;
  assign new_n2284_ = ~new_n2239_;
  assign new_n2285_ = ~new_n2239_ | ~new_n1956_;
  assign new_n2286_ = ~new_n2238_ | ~new_n1957_;
  assign po068 = new_n2241_;
  assign new_n2288_ = ~new_n2241_;
  assign new_n2289_ = ~new_n2242_ | ~new_n2184_;
  assign new_n2290_ = ~new_n2243_ | ~new_n2185_;
  assign new_n2291_ = ~new_n1983_ | ~new_n2229_;
  assign po069 = new_n2244_;
  assign new_n2293_ = ~new_n2244_;
  assign new_n2294_ = new_n729_ | new_n911_ | new_n2221_ | new_n2225_;
  assign new_n2295_ = new_n730_ | new_n910_ | new_n2214_ | new_n2218_;
  assign new_n2296_ = new_n737_ | new_n919_ | new_n2156_ | new_n2217_;
  assign new_n2297_ = new_n738_ | new_n918_ | new_n2158_ | new_n2224_;
  assign new_n2298_ = new_n739_ | new_n925_ | new_n2219_ | new_n2223_;
  assign new_n2299_ = new_n740_ | new_n924_ | new_n2212_ | new_n2216_;
  assign new_n2300_ = new_n741_ | new_n927_ | new_n2213_ | new_n2215_;
  assign new_n2301_ = new_n742_ | new_n926_ | new_n2220_ | new_n2222_;
  assign po072 = new_n2245_ & new_n747_;
  assign po073 = new_n2246_ & new_n749_;
  assign new_n2304_ = new_n941_ | new_n1410_ | new_n2196_;
  assign po100 = ~new_n2253_;
  assign po095 = ~new_n2254_;
  assign po081 = new_n766_ | new_n958_ | new_n2152_ | new_n2204_;
  assign po077 = new_n767_ | new_n959_ | new_n2155_ | new_n2209_;
  assign new_n2309_ = new_n960_ | new_n1413_ | new_n2197_;
  assign po078 = new_n777_ | new_n964_ | new_n2198_ | new_n2201_;
  assign po074 = new_n778_ | new_n965_ | new_n2206_ | new_n2205_;
  assign po079 = new_n782_ | new_n954_ | new_n2199_ | new_n2202_;
  assign po075 = new_n783_ | new_n955_ | new_n2210_ | new_n2207_;
  assign po076 = new_n784_ | new_n956_ | new_n2211_ | new_n2208_;
  assign po080 = new_n785_ | new_n957_ | new_n2200_ | new_n2203_;
  assign new_n2316_ = new_n2278_ & new_n501_;
  assign new_n2317_ = new_n2277_ & new_n501_;
  assign new_n2318_ = new_n502_ & new_n2304_ & new_n504_;
  assign new_n2319_ = new_n502_ & new_n2309_ & new_n314_;
  assign new_n2320_ = new_n508_ & new_n2309_ & new_n316_;
  assign new_n2321_ = new_n508_ & new_n2304_ & new_n506_;
  assign new_n2322_ = new_n524_ & new_n2304_ & new_n526_;
  assign new_n2323_ = new_n524_ & new_n2309_ & new_n335_;
  assign new_n2324_ = new_n528_ & new_n2304_ & new_n530_;
  assign new_n2325_ = new_n528_ & new_n2309_ & new_n339_;
  assign new_n2326_ = new_n2102_ & new_n2045_ & new_n2293_ & pi155 & new_n2288_;
  assign new_n2327_ = ~new_n1792_ | ~new_n2271_;
  assign new_n2328_ = ~new_n2273_;
  assign new_n2329_ = new_n2291_ & new_n2229_;
  assign new_n2330_ = ~new_n2277_;
  assign new_n2331_ = ~new_n2289_ | ~new_n1802_;
  assign new_n2332_ = ~new_n2290_ | ~new_n1803_;
  assign new_n2333_ = ~new_n2278_;
  assign new_n2334_ = ~new_n2279_;
  assign new_n2335_ = ~new_n2280_;
  assign new_n2336_ = ~new_n2279_ | ~new_n1848_;
  assign new_n2337_ = ~new_n2280_ | ~new_n1849_;
  assign new_n2338_ = ~new_n1866_ | ~new_n2284_;
  assign new_n2339_ = ~new_n1867_ | ~new_n2283_;
  assign new_n2340_ = ~new_n2273_ | ~new_n1490_;
  assign new_n2341_ = ~new_n2289_;
  assign new_n2342_ = ~new_n2290_;
  assign new_n2343_ = new_n1983_ & new_n2291_;
  assign new_n2344_ = new_n727_ | new_n908_ | new_n2267_ | new_n2268_;
  assign new_n2345_ = new_n728_ | new_n909_ | new_n2269_ | new_n2270_;
  assign po082 = new_n2294_ & new_n746_;
  assign po083 = new_n2297_ & new_n747_;
  assign po084 = new_n2298_ & new_n747_;
  assign po085 = new_n2301_ & new_n747_;
  assign po087 = new_n2296_ & new_n749_;
  assign po088 = new_n2299_ & new_n749_;
  assign po089 = new_n2300_ & new_n749_;
  assign po086 = new_n2295_ & new_n750_;
  assign new_n2354_ = new_n2266_ | new_n753_ | new_n1245_ | new_n1992_;
  assign new_n2355_ = new_n934_ | new_n1243_ | new_n2258_;
  assign new_n2356_ = new_n936_ | new_n1242_ | new_n2259_;
  assign po094 = ~new_n2304_;
  assign new_n2358_ = new_n942_ | new_n1525_ | new_n2260_;
  assign new_n2359_ = new_n943_ | new_n1414_ | new_n2261_;
  assign po071 = new_n2275_ & new_n2274_ & new_n2230_ & new_n2169_ & new_n2115_ & new_n2114_ & new_n2112_ & new_n1900_ & new_n2091_;
  assign po099 = ~new_n2309_;
  assign po105 = new_n775_ | new_n951_ | new_n2265_ | new_n2264_;
  assign po108 = new_n776_ | new_n950_ | new_n2262_ | new_n2263_;
  assign po070 = new_n2282_ & new_n2281_ & new_n2237_ & new_n2176_ & new_n2125_ & new_n2136_ & new_n2132_ & new_n2103_ & new_n2133_;
  assign new_n2365_ = new_n493_ & new_n2330_ & new_n499_;
  assign new_n2366_ = new_n495_ & new_n2333_ & new_n500_;
  assign new_n2367_ = new_n502_ & new_n2355_ & new_n504_;
  assign new_n2368_ = new_n502_ & new_n2356_ & new_n504_;
  assign new_n2369_ = new_n502_ & new_n2358_ & new_n314_;
  assign new_n2370_ = new_n502_ & new_n2359_ & new_n314_;
  assign new_n2371_ = new_n508_ & new_n2358_ & new_n316_;
  assign new_n2372_ = new_n508_ & new_n2359_ & new_n316_;
  assign new_n2373_ = new_n508_ & new_n2355_ & new_n506_;
  assign new_n2374_ = new_n508_ & new_n2356_ & new_n506_;
  assign new_n2375_ = new_n524_ & new_n2356_ & new_n526_;
  assign new_n2376_ = new_n524_ & new_n2355_ & new_n526_;
  assign new_n2377_ = new_n524_ & new_n2358_ & new_n335_;
  assign new_n2378_ = new_n524_ & new_n2359_ & new_n335_;
  assign new_n2379_ = new_n528_ & new_n2356_ & new_n530_;
  assign new_n2380_ = new_n528_ & new_n2355_ & new_n530_;
  assign new_n2381_ = new_n528_ & new_n2358_ & new_n339_;
  assign new_n2382_ = new_n528_ & new_n2359_ & new_n339_;
  assign new_n2383_ = ~new_n2327_ | ~new_n2272_;
  assign po091 = new_n2343_ | new_n2329_;
  assign new_n2385_ = ~new_n1624_ | ~new_n2341_;
  assign new_n2386_ = ~new_n1626_ | ~new_n2342_;
  assign new_n2387_ = ~new_n1684_ | ~new_n2334_;
  assign new_n2388_ = ~new_n1685_ | ~new_n2335_;
  assign new_n2389_ = ~new_n2338_ | ~new_n2285_;
  assign new_n2390_ = ~new_n2339_ | ~new_n2286_;
  assign new_n2391_ = ~new_n1324_ | ~new_n2328_;
  assign po096 = pi098 & new_n379_ & new_n2326_;
  assign new_n2393_ = new_n731_ | new_n913_ | new_n2324_ | new_n2325_;
  assign new_n2394_ = new_n732_ | new_n912_ | new_n2322_ | new_n2323_;
  assign po109 = new_n2345_ & new_n746_;
  assign po113 = new_n2344_ & new_n750_;
  assign po090 = new_n752_ & new_n2354_;
  assign po092 = ~new_n2355_;
  assign po093 = ~new_n2356_;
  assign po097 = ~new_n2358_;
  assign po098 = ~new_n2359_;
  assign po107 = new_n756_ | new_n948_ | new_n2318_ | new_n2319_;
  assign po104 = new_n757_ | new_n949_ | new_n2321_ | new_n2320_;
  assign new_n2404_ = ~new_n2383_;
  assign new_n2405_ = ~new_n2385_ | ~new_n2331_;
  assign new_n2406_ = ~new_n2386_ | ~new_n2332_;
  assign new_n2407_ = ~new_n2387_ | ~new_n2336_;
  assign new_n2408_ = ~new_n2388_ | ~new_n2337_;
  assign new_n2409_ = ~new_n2389_;
  assign new_n2410_ = ~new_n2390_;
  assign new_n2411_ = ~new_n2389_ | ~new_n1868_;
  assign new_n2412_ = ~new_n2390_ | ~new_n1869_;
  assign new_n2413_ = ~new_n2383_ | ~new_n1489_;
  assign new_n2414_ = ~new_n2391_ | ~new_n2340_;
  assign new_n2415_ = new_n733_ | new_n914_ | new_n2375_ | new_n2378_;
  assign new_n2416_ = new_n734_ | new_n915_ | new_n2379_ | new_n2382_;
  assign new_n2417_ = new_n735_ | new_n917_ | new_n2380_ | new_n2381_;
  assign new_n2418_ = new_n736_ | new_n916_ | new_n2376_ | new_n2377_;
  assign po110 = new_n2393_ & new_n746_;
  assign po114 = new_n2394_ & new_n750_;
  assign po101 = new_n754_ | new_n946_ | new_n2367_ | new_n2369_;
  assign po102 = new_n755_ | new_n947_ | new_n2373_ | new_n2371_;
  assign po106 = new_n773_ | new_n962_ | new_n2368_ | new_n2370_;
  assign po103 = new_n774_ | new_n963_ | new_n2374_ | new_n2372_;
  assign new_n2425_ = ~new_n2414_ | ~new_n1779_;
  assign new_n2426_ = ~new_n2405_;
  assign new_n2427_ = ~new_n2406_;
  assign new_n2428_ = ~new_n2406_ | ~new_n1810_;
  assign new_n2429_ = ~new_n2405_ | ~new_n1811_;
  assign new_n2430_ = ~new_n2408_ | ~new_n1819_;
  assign new_n2431_ = ~new_n2407_ | ~new_n1821_;
  assign new_n2432_ = ~new_n2407_;
  assign new_n2433_ = ~new_n2408_;
  assign new_n2434_ = ~new_n1718_ | ~new_n2409_;
  assign new_n2435_ = ~new_n1719_ | ~new_n2410_;
  assign new_n2436_ = ~new_n1323_ | ~new_n2404_;
  assign new_n2437_ = ~new_n2414_;
  assign po111 = new_n2416_ & new_n746_;
  assign po112 = new_n2417_ & new_n746_;
  assign po115 = new_n2415_ & new_n750_;
  assign po116 = new_n2418_ & new_n750_;
  assign new_n2442_ = ~new_n1598_ | ~new_n2437_;
  assign new_n2443_ = ~new_n1640_ | ~new_n2427_;
  assign new_n2444_ = ~new_n1641_ | ~new_n2426_;
  assign new_n2445_ = ~new_n1653_ | ~new_n2433_;
  assign new_n2446_ = ~new_n1656_ | ~new_n2432_;
  assign new_n2447_ = ~new_n2434_ | ~new_n2411_;
  assign new_n2448_ = ~new_n2435_ | ~new_n2412_;
  assign new_n2449_ = ~new_n2436_ | ~new_n2413_;
  assign new_n2450_ = ~new_n2442_ | ~new_n2425_;
  assign new_n2451_ = ~new_n2449_ | ~new_n1780_;
  assign new_n2452_ = ~new_n2443_ | ~new_n2428_;
  assign new_n2453_ = ~new_n2444_ | ~new_n2429_;
  assign new_n2454_ = ~new_n2445_ | ~new_n2430_;
  assign new_n2455_ = ~new_n2446_ | ~new_n2431_;
  assign new_n2456_ = ~new_n2448_ | ~new_n1853_;
  assign new_n2457_ = ~new_n2447_ | ~new_n1854_;
  assign new_n2458_ = ~new_n2447_;
  assign new_n2459_ = ~new_n2448_;
  assign new_n2460_ = ~new_n2449_;
  assign new_n2461_ = ~new_n2450_;
  assign new_n2462_ = ~new_n1599_ | ~new_n2460_;
  assign new_n2463_ = ~new_n2450_ | ~new_n1796_;
  assign new_n2464_ = ~new_n2452_;
  assign new_n2465_ = ~new_n2453_;
  assign new_n2466_ = ~new_n2454_;
  assign new_n2467_ = ~new_n2455_;
  assign new_n2468_ = ~new_n2455_ | ~new_n1836_;
  assign new_n2469_ = ~new_n2454_ | ~new_n1837_;
  assign new_n2470_ = ~new_n1695_ | ~new_n2459_;
  assign new_n2471_ = ~new_n1698_ | ~new_n2458_;
  assign new_n2472_ = ~new_n2453_ | ~new_n1507_;
  assign new_n2473_ = ~new_n2452_ | ~new_n1508_;
  assign new_n2474_ = ~new_n2462_ | ~new_n2451_;
  assign new_n2475_ = ~new_n1621_ | ~new_n2461_;
  assign new_n2476_ = ~new_n1670_ | ~new_n2467_;
  assign new_n2477_ = ~new_n1671_ | ~new_n2466_;
  assign new_n2478_ = ~new_n2470_ | ~new_n2456_;
  assign new_n2479_ = ~new_n2471_ | ~new_n2457_;
  assign new_n2480_ = ~new_n1361_ | ~new_n2465_;
  assign new_n2481_ = ~new_n1362_ | ~new_n2464_;
  assign new_n2482_ = ~new_n2474_;
  assign new_n2483_ = ~new_n2474_ | ~new_n1795_;
  assign new_n2484_ = ~new_n2475_ | ~new_n2463_;
  assign new_n2485_ = ~new_n2476_ | ~new_n2468_;
  assign new_n2486_ = ~new_n2477_ | ~new_n2469_;
  assign new_n2487_ = ~new_n2479_ | ~new_n1840_;
  assign new_n2488_ = ~new_n2478_ | ~new_n1841_;
  assign new_n2489_ = ~new_n2478_;
  assign new_n2490_ = ~new_n2479_;
  assign new_n2491_ = ~new_n2480_ | ~new_n2472_;
  assign new_n2492_ = ~new_n2481_ | ~new_n2473_;
  assign new_n2493_ = ~new_n2484_ | ~new_n1787_;
  assign new_n2494_ = ~new_n1620_ | ~new_n2482_;
  assign new_n2495_ = ~new_n2484_;
  assign new_n2496_ = ~new_n2486_ | ~new_n1824_;
  assign new_n2497_ = ~new_n2485_ | ~new_n1825_;
  assign new_n2498_ = ~new_n2485_;
  assign new_n2499_ = ~new_n2486_;
  assign new_n2500_ = ~new_n1673_ | ~new_n2490_;
  assign new_n2501_ = ~new_n1674_ | ~new_n2489_;
  assign new_n2502_ = ~new_n2492_ | ~new_n1502_;
  assign new_n2503_ = ~new_n2491_ | ~new_n1503_;
  assign new_n2504_ = ~new_n2491_;
  assign new_n2505_ = ~new_n2492_;
  assign new_n2506_ = ~new_n1612_ | ~new_n2495_;
  assign new_n2507_ = ~new_n2494_ | ~new_n2483_;
  assign new_n2508_ = ~new_n1661_ | ~new_n2499_;
  assign new_n2509_ = ~new_n1662_ | ~new_n2498_;
  assign new_n2510_ = ~new_n2500_ | ~new_n2487_;
  assign new_n2511_ = ~new_n2501_ | ~new_n2488_;
  assign new_n2512_ = ~new_n1351_ | ~new_n2505_;
  assign new_n2513_ = ~new_n1352_ | ~new_n2504_;
  assign new_n2514_ = ~new_n2507_ | ~new_n1786_;
  assign new_n2515_ = ~new_n2506_ | ~new_n2493_;
  assign new_n2516_ = ~new_n2507_;
  assign new_n2517_ = ~new_n2508_ | ~new_n2496_;
  assign new_n2518_ = ~new_n2509_ | ~new_n2497_;
  assign new_n2519_ = ~new_n2510_;
  assign new_n2520_ = ~new_n2511_;
  assign new_n2521_ = ~new_n2510_ | ~new_n1856_;
  assign new_n2522_ = ~new_n2511_ | ~new_n1857_;
  assign new_n2523_ = ~new_n2512_ | ~new_n2502_;
  assign new_n2524_ = ~new_n2513_ | ~new_n2503_;
  assign new_n2525_ = new_n331_ & new_n2524_ & new_n1916_;
  assign new_n2526_ = new_n331_ & new_n2523_ & new_n1797_;
  assign new_n2527_ = pi161 & new_n2523_ & new_n2093_;
  assign new_n2528_ = pi161 & new_n2524_ & new_n2040_;
  assign new_n2529_ = new_n340_ & new_n2518_ & new_n1941_;
  assign new_n2530_ = new_n340_ & new_n2517_ & new_n1843_;
  assign new_n2531_ = pi156 & new_n2517_ & new_n2076_;
  assign new_n2532_ = pi156 & new_n2518_ & new_n2019_;
  assign new_n2533_ = ~new_n1611_ | ~new_n2516_;
  assign new_n2534_ = ~new_n2515_;
  assign new_n2535_ = ~new_n2515_ | ~new_n1616_;
  assign new_n2536_ = ~new_n1705_ | ~new_n2519_;
  assign new_n2537_ = ~new_n1706_ | ~new_n2520_;
  assign new_n2538_ = new_n2527_ | new_n2528_ | new_n2525_ | new_n2526_;
  assign new_n2539_ = new_n2531_ | new_n2532_ | new_n2529_ | new_n2530_;
  assign new_n2540_ = ~new_n2533_ | ~new_n2514_;
  assign new_n2541_ = ~new_n1538_ | ~new_n2534_;
  assign new_n2542_ = ~new_n2536_ | ~new_n2521_;
  assign new_n2543_ = ~new_n2537_ | ~new_n2522_;
  assign new_n2544_ = ~new_n2538_;
  assign new_n2545_ = ~new_n2539_;
  assign new_n2546_ = ~new_n2540_;
  assign new_n2547_ = ~new_n2540_ | ~new_n1615_;
  assign new_n2548_ = ~new_n2541_ | ~new_n2535_;
  assign new_n2549_ = ~new_n2542_;
  assign new_n2550_ = ~new_n2543_;
  assign new_n2551_ = ~new_n2542_ | ~new_n1864_;
  assign new_n2552_ = ~new_n2543_ | ~new_n1865_;
  assign new_n2553_ = pi161 & new_n2548_;
  assign new_n2554_ = ~new_n1537_ | ~new_n2546_;
  assign new_n2555_ = ~new_n1715_ | ~new_n2549_;
  assign new_n2556_ = ~new_n1716_ | ~new_n2550_;
  assign new_n2557_ = ~new_n2554_ | ~new_n2547_;
  assign new_n2558_ = ~new_n2555_ | ~new_n2551_;
  assign new_n2559_ = ~new_n2556_ | ~new_n2552_;
  assign new_n2560_ = pi156 & new_n2559_;
  assign new_n2561_ = ~new_n2557_;
  assign new_n2562_ = ~new_n2558_;
  assign new_n2563_ = new_n2561_ & new_n331_;
  assign new_n2564_ = new_n2562_ & new_n340_;
  assign new_n2565_ = new_n2563_ | new_n2553_;
  assign new_n2566_ = new_n2564_ | new_n2560_;
  assign new_n2567_ = ~new_n2565_ | ~new_n2544_;
  assign new_n2568_ = ~new_n2565_;
  assign new_n2569_ = ~new_n2566_ | ~new_n2545_;
  assign new_n2570_ = ~new_n2566_;
  assign new_n2571_ = ~new_n2538_ | ~new_n2568_;
  assign new_n2572_ = ~new_n2539_ | ~new_n2570_;
  assign new_n2573_ = ~new_n2567_ | ~new_n2571_;
  assign new_n2574_ = ~new_n2569_ | ~new_n2572_;
  assign new_n2575_ = new_n493_ & new_n2573_ & new_n309_;
  assign new_n2576_ = new_n495_ & new_n2574_ & new_n310_;
  assign new_n2577_ = ~new_n2573_;
  assign new_n2578_ = ~new_n2574_;
  assign po117 = new_n492_ | new_n937_ | new_n2365_ | new_n2575_;
  assign po118 = new_n494_ | new_n939_ | new_n2366_ | new_n2576_;
  assign new_n2581_ = new_n2577_ & new_n311_;
  assign new_n2582_ = new_n2578_ & new_n311_;
  assign new_n2583_ = new_n2316_ | new_n2582_;
  assign new_n2584_ = new_n2317_ | new_n2581_;
  assign new_n2585_ = new_n2583_ & new_n496_;
  assign new_n2586_ = new_n2583_ & new_n496_;
  assign new_n2587_ = new_n2584_ & new_n496_;
  assign new_n2588_ = new_n2584_ & new_n496_;
  assign new_n2589_ = new_n2586_ | new_n758_;
  assign new_n2590_ = new_n2585_ | new_n759_;
  assign new_n2591_ = new_n2588_ | new_n760_;
  assign new_n2592_ = new_n2587_ | new_n761_;
  assign new_n2593_ = new_n503_ & new_n2591_ & new_n505_;
  assign new_n2594_ = new_n503_ & new_n2589_ & new_n315_;
  assign new_n2595_ = new_n509_ & new_n2589_ & new_n317_;
  assign new_n2596_ = new_n509_ & new_n2591_ & new_n507_;
  assign new_n2597_ = new_n523_ & new_n2592_ & new_n525_;
  assign new_n2598_ = new_n523_ & new_n2590_ & new_n334_;
  assign new_n2599_ = new_n527_ & new_n2592_ & new_n529_;
  assign new_n2600_ = new_n527_ & new_n2590_ & new_n338_;
  assign new_n2601_ = new_n725_ | new_n923_ | new_n2599_ | new_n2600_;
  assign new_n2602_ = new_n726_ | new_n922_ | new_n2597_ | new_n2598_;
  assign po119 = new_n768_ | new_n971_ | new_n2596_ | new_n2595_;
  assign po120 = new_n769_ | new_n970_ | new_n2593_ | new_n2594_;
  assign new_n2605_ = new_n2601_ & new_n747_;
  assign new_n2606_ = new_n2602_ & new_n749_;
  assign po121 = ~new_n2605_;
  assign po122 = ~new_n2606_;
endmodule


