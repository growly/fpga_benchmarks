// Benchmark "i9" written by ABC on Thu Mar 19 13:02:36 2020

module i9 ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47,
    pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71,
    pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81, pi82, pi83,
    pi84, pi85, pi86, pi87,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47,
    po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45,
    pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57,
    pi58, pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69,
    pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81,
    pi82, pi83, pi84, pi85, pi86, pi87;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46,
    po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58,
    po59, po60, po61, po62;
  wire new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_,
    new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_,
    new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_,
    new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_,
    new_n176_, new_n178_, new_n180_, new_n182_, new_n184_, new_n186_,
    new_n188_, new_n190_, new_n192_, new_n194_, new_n196_, new_n198_,
    new_n200_, new_n202_, new_n204_, new_n206_, new_n208_, new_n210_,
    new_n212_, new_n214_, new_n216_, new_n218_, new_n220_, new_n222_,
    new_n224_, new_n226_, new_n228_, new_n230_, new_n232_, new_n234_,
    new_n236_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_;
  assign new_n152_ = pi02 & pi00 & pi01;
  assign new_n153_ = pi03 & pi01;
  assign new_n154_ = pi03 & pi02;
  assign new_n155_ = ~pi04;
  assign new_n156_ = ~pi05;
  assign new_n157_ = ~pi03;
  assign new_n158_ = new_n156_ & new_n157_ & new_n155_;
  assign new_n159_ = ~pi02;
  assign new_n160_ = ~pi06;
  assign new_n161_ = new_n160_ & new_n159_ & pi01 & new_n157_ & new_n156_;
  assign new_n162_ = pi07 & new_n157_ & new_n155_;
  assign new_n163_ = pi08 & new_n157_ & pi01;
  assign new_n164_ = ~pi00;
  assign new_n165_ = new_n164_ & pi01 & new_n157_ & pi02;
  assign new_n166_ = ~pi01;
  assign new_n167_ = new_n160_ & pi02 & pi04 & new_n166_ & new_n157_ & new_n156_;
  assign new_n168_ = pi08 & new_n166_ & new_n157_ & pi02;
  assign new_n169_ = new_n156_ & new_n166_ & new_n160_ & new_n159_;
  assign new_n170_ = new_n159_ & pi07 & new_n166_;
  assign new_n171_ = new_n159_ & pi03 & new_n166_;
  assign new_n172_ = new_n168_ | new_n165_ | new_n167_ | new_n163_ | new_n158_ | new_n161_ | new_n162_ | new_n153_ | new_n152_ | new_n169_ | new_n154_ | new_n171_ | new_n170_;
  assign new_n173_ = new_n171_ | new_n170_ | new_n169_ | new_n165_ | new_n168_ | new_n167_;
  assign new_n174_ = new_n171_ | new_n170_ | new_n169_ | new_n158_ | new_n161_ | new_n163_ | new_n162_;
  assign new_n175_ = ~new_n172_;
  assign new_n176_ = new_n172_ & new_n484_ & pi09 & new_n485_;
  assign po00 = new_n262_ | new_n293_ | new_n238_ | new_n175_ | new_n176_;
  assign new_n178_ = new_n172_ & new_n484_ & pi10 & new_n485_;
  assign po01 = new_n263_ | new_n294_ | new_n239_ | new_n175_ | new_n178_;
  assign new_n180_ = new_n172_ & new_n484_ & pi11 & new_n485_;
  assign po02 = new_n264_ | new_n295_ | new_n240_ | new_n175_ | new_n180_;
  assign new_n182_ = new_n172_ & new_n484_ & pi12 & new_n485_;
  assign po03 = new_n265_ | new_n296_ | new_n241_ | new_n175_ | new_n182_;
  assign new_n184_ = new_n172_ & new_n484_ & pi13 & new_n485_;
  assign po04 = new_n266_ | new_n297_ | new_n242_ | new_n175_ | new_n184_;
  assign new_n186_ = new_n172_ & new_n484_ & pi14 & new_n485_;
  assign po05 = new_n267_ | new_n298_ | new_n243_ | new_n175_ | new_n186_;
  assign new_n188_ = new_n172_ & new_n484_ & pi15 & new_n485_;
  assign po06 = new_n268_ | new_n299_ | new_n244_ | new_n175_ | new_n188_;
  assign new_n190_ = new_n172_ & new_n484_ & pi16 & new_n485_;
  assign po07 = new_n269_ | new_n300_ | new_n245_ | new_n175_ | new_n190_;
  assign new_n192_ = new_n172_ & new_n484_ & pi17 & new_n485_;
  assign po08 = new_n270_ | new_n301_ | new_n246_ | new_n175_ | new_n192_;
  assign new_n194_ = new_n172_ & new_n484_ & pi18 & new_n485_;
  assign po09 = new_n271_ | new_n302_ | new_n247_ | new_n175_ | new_n194_;
  assign new_n196_ = new_n172_ & new_n484_ & pi19 & new_n485_;
  assign po10 = new_n272_ | new_n303_ | new_n248_ | new_n175_ | new_n196_;
  assign new_n198_ = new_n172_ & new_n484_ & pi20 & new_n485_;
  assign po11 = new_n273_ | new_n304_ | new_n249_ | new_n175_ | new_n198_;
  assign new_n200_ = new_n172_ & new_n484_ & pi21 & new_n485_;
  assign po12 = new_n274_ | new_n305_ | new_n250_ | new_n175_ | new_n200_;
  assign new_n202_ = new_n172_ & new_n484_ & pi22 & new_n485_;
  assign po13 = new_n275_ | new_n306_ | new_n251_ | new_n175_ | new_n202_;
  assign new_n204_ = new_n172_ & new_n484_ & pi23 & new_n485_;
  assign po14 = new_n276_ | new_n307_ | new_n252_ | new_n175_ | new_n204_;
  assign new_n206_ = new_n172_ & new_n484_ & pi24 & new_n485_;
  assign po15 = new_n277_ | new_n308_ | new_n253_ | new_n175_ | new_n206_;
  assign new_n208_ = new_n172_ & new_n484_ & pi25 & new_n485_;
  assign po16 = new_n278_ | new_n309_ | new_n254_ | new_n175_ | new_n208_;
  assign new_n210_ = new_n172_ & new_n484_ & pi26 & new_n485_;
  assign po17 = new_n279_ | new_n310_ | new_n255_ | new_n175_ | new_n210_;
  assign new_n212_ = new_n172_ & new_n484_ & pi27 & new_n485_;
  assign po18 = new_n280_ | new_n311_ | new_n256_ | new_n175_ | new_n212_;
  assign new_n214_ = new_n172_ & new_n484_ & pi28 & new_n485_;
  assign po19 = new_n281_ | new_n312_ | new_n257_ | new_n175_ | new_n214_;
  assign new_n216_ = new_n172_ & new_n484_ & pi29 & new_n485_;
  assign po20 = new_n282_ | new_n313_ | new_n258_ | new_n175_ | new_n216_;
  assign new_n218_ = new_n172_ & new_n484_ & pi30 & new_n485_;
  assign po21 = new_n283_ | new_n314_ | new_n259_ | new_n175_ | new_n218_;
  assign new_n220_ = new_n172_ & new_n484_ & pi31 & new_n485_;
  assign po22 = new_n284_ | new_n315_ | new_n260_ | new_n175_ | new_n220_;
  assign new_n222_ = new_n172_ & new_n484_ & pi32 & new_n485_;
  assign po23 = new_n285_ | new_n316_ | new_n261_ | new_n175_ | new_n222_;
  assign new_n224_ = new_n172_ & new_n484_ & pi33 & new_n485_;
  assign po24 = new_n286_ | new_n317_ | new_n487_ | new_n175_ | new_n224_;
  assign new_n226_ = new_n172_ & new_n484_ & pi34 & new_n485_;
  assign po25 = new_n287_ | new_n318_ | new_n487_ | new_n175_ | new_n226_;
  assign new_n228_ = new_n172_ & new_n484_ & pi35 & new_n485_;
  assign po26 = new_n288_ | new_n319_ | new_n487_ | new_n175_ | new_n228_;
  assign new_n230_ = new_n172_ & new_n484_ & pi36 & new_n485_;
  assign po27 = new_n289_ | new_n320_ | new_n487_ | new_n175_ | new_n230_;
  assign new_n232_ = new_n172_ & new_n484_ & pi37 & new_n485_;
  assign po28 = new_n290_ | new_n321_ | new_n487_ | new_n175_ | new_n232_;
  assign new_n234_ = new_n172_ & new_n484_ & pi38 & new_n485_;
  assign po29 = new_n291_ | new_n322_ | new_n487_ | new_n175_ | new_n234_;
  assign new_n236_ = new_n172_ & new_n484_ & pi39 & new_n485_;
  assign po30 = new_n292_ | new_n323_ | new_n487_ | new_n175_ | new_n236_;
  assign new_n238_ = new_n487_ & pi17;
  assign new_n239_ = new_n487_ & pi18;
  assign new_n240_ = new_n487_ & pi19;
  assign new_n241_ = new_n487_ & pi20;
  assign new_n242_ = new_n487_ & pi21;
  assign new_n243_ = new_n487_ & pi22;
  assign new_n244_ = new_n487_ & pi23;
  assign new_n245_ = new_n487_ & pi24;
  assign new_n246_ = new_n487_ & pi25;
  assign new_n247_ = new_n487_ & pi26;
  assign new_n248_ = new_n487_ & pi27;
  assign new_n249_ = new_n487_ & pi28;
  assign new_n250_ = new_n487_ & pi29;
  assign new_n251_ = new_n487_ & pi30;
  assign new_n252_ = new_n487_ & pi31;
  assign new_n253_ = new_n487_ & pi32;
  assign new_n254_ = new_n487_ & pi33;
  assign new_n255_ = new_n487_ & pi34;
  assign new_n256_ = new_n487_ & pi35;
  assign new_n257_ = new_n487_ & pi36;
  assign new_n258_ = new_n487_ & pi37;
  assign new_n259_ = new_n487_ & pi38;
  assign new_n260_ = new_n487_ & pi39;
  assign new_n261_ = new_n487_ & pi40;
  assign new_n262_ = new_n172_ & new_n173_ & pi20 & new_n488_;
  assign new_n263_ = new_n172_ & new_n173_ & pi21 & new_n488_;
  assign new_n264_ = new_n172_ & new_n173_ & pi22 & new_n488_;
  assign new_n265_ = new_n172_ & new_n173_ & pi23 & new_n488_;
  assign new_n266_ = new_n172_ & new_n173_ & pi24 & new_n488_;
  assign new_n267_ = new_n172_ & new_n173_ & pi25 & new_n488_;
  assign new_n268_ = new_n172_ & new_n173_ & pi26 & new_n488_;
  assign new_n269_ = new_n172_ & new_n173_ & pi27 & new_n488_;
  assign new_n270_ = new_n172_ & new_n173_ & pi28 & new_n488_;
  assign new_n271_ = new_n172_ & new_n173_ & pi29 & new_n488_;
  assign new_n272_ = new_n172_ & new_n173_ & pi30 & new_n488_;
  assign new_n273_ = new_n172_ & new_n173_ & pi31 & new_n488_;
  assign new_n274_ = new_n172_ & new_n173_ & pi32 & new_n488_;
  assign new_n275_ = new_n172_ & new_n173_ & pi33 & new_n488_;
  assign new_n276_ = new_n172_ & new_n173_ & pi34 & new_n488_;
  assign new_n277_ = new_n172_ & new_n173_ & pi35 & new_n488_;
  assign new_n278_ = new_n172_ & new_n173_ & pi36 & new_n488_;
  assign new_n279_ = new_n172_ & new_n173_ & pi37 & new_n488_;
  assign new_n280_ = new_n172_ & new_n173_ & pi38 & new_n488_;
  assign new_n281_ = new_n172_ & new_n173_ & pi39 & new_n488_;
  assign new_n282_ = new_n172_ & new_n173_ & pi41 & new_n488_;
  assign new_n283_ = new_n172_ & new_n173_ & pi42 & new_n488_;
  assign new_n284_ = new_n172_ & new_n173_ & pi43 & new_n488_;
  assign new_n285_ = new_n172_ & new_n173_ & pi44 & new_n488_;
  assign new_n286_ = new_n172_ & new_n173_ & pi45 & new_n488_;
  assign new_n287_ = new_n172_ & new_n173_ & pi46 & new_n488_;
  assign new_n288_ = new_n172_ & new_n173_ & pi47 & new_n488_;
  assign new_n289_ = new_n172_ & new_n173_ & pi48 & new_n488_;
  assign new_n290_ = new_n172_ & new_n173_ & pi49 & new_n488_;
  assign new_n291_ = new_n172_ & new_n173_ & pi50 & new_n488_;
  assign new_n292_ = new_n172_ & new_n173_ & pi51 & new_n488_;
  assign new_n293_ = new_n172_ & new_n173_ & pi24 & new_n174_;
  assign new_n294_ = new_n172_ & new_n173_ & pi25 & new_n174_;
  assign new_n295_ = new_n172_ & new_n173_ & pi26 & new_n174_;
  assign new_n296_ = new_n172_ & new_n173_ & pi27 & new_n174_;
  assign new_n297_ = new_n172_ & new_n173_ & pi28 & new_n174_;
  assign new_n298_ = new_n172_ & new_n173_ & pi29 & new_n174_;
  assign new_n299_ = new_n172_ & new_n173_ & pi30 & new_n174_;
  assign new_n300_ = new_n172_ & new_n173_ & pi31 & new_n174_;
  assign new_n301_ = new_n172_ & new_n173_ & pi32 & new_n174_;
  assign new_n302_ = new_n172_ & new_n173_ & pi33 & new_n174_;
  assign new_n303_ = new_n172_ & new_n173_ & pi34 & new_n174_;
  assign new_n304_ = new_n172_ & new_n173_ & pi35 & new_n174_;
  assign new_n305_ = new_n172_ & new_n173_ & pi36 & new_n174_;
  assign new_n306_ = new_n172_ & new_n173_ & pi37 & new_n174_;
  assign new_n307_ = new_n172_ & new_n173_ & pi38 & new_n174_;
  assign new_n308_ = new_n172_ & new_n173_ & pi39 & new_n174_;
  assign new_n309_ = new_n172_ & new_n173_ & pi52 & new_n174_;
  assign new_n310_ = new_n172_ & new_n173_ & pi53 & new_n174_;
  assign new_n311_ = new_n172_ & new_n173_ & pi54 & new_n174_;
  assign new_n312_ = new_n172_ & new_n173_ & pi55 & new_n174_;
  assign new_n313_ = new_n172_ & new_n173_ & pi56 & new_n174_;
  assign new_n314_ = new_n172_ & new_n173_ & pi57 & new_n174_;
  assign new_n315_ = new_n172_ & new_n173_ & pi58 & new_n174_;
  assign new_n316_ = new_n172_ & new_n173_ & pi59 & new_n174_;
  assign new_n317_ = new_n172_ & new_n173_ & pi60 & new_n174_;
  assign new_n318_ = new_n172_ & new_n173_ & pi61 & new_n174_;
  assign new_n319_ = new_n172_ & new_n173_ & pi62 & new_n174_;
  assign new_n320_ = new_n172_ & new_n173_ & pi63 & new_n174_;
  assign new_n321_ = new_n172_ & new_n173_ & pi64 & new_n174_;
  assign new_n322_ = new_n172_ & new_n173_ & pi65 & new_n174_;
  assign new_n323_ = new_n172_ & new_n173_ & pi66 & new_n174_;
  assign po31 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n372_ | new_n404_ | new_n436_ | new_n468_;
  assign po32 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n373_ | new_n405_ | new_n437_ | new_n469_;
  assign po33 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n374_ | new_n406_ | new_n438_ | new_n470_;
  assign po34 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n375_ | new_n407_ | new_n439_ | new_n471_;
  assign po35 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n376_ | new_n408_ | new_n440_ | new_n472_;
  assign po36 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n377_ | new_n409_ | new_n441_ | new_n473_;
  assign po37 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n378_ | new_n410_ | new_n442_ | new_n474_;
  assign po38 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n379_ | new_n411_ | new_n443_ | new_n475_;
  assign po39 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n380_ | new_n412_ | new_n444_ | new_n476_;
  assign po40 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n381_ | new_n413_ | new_n445_ | new_n477_;
  assign po41 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n382_ | new_n414_ | new_n446_ | new_n478_;
  assign po42 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n383_ | new_n415_ | new_n447_ | new_n479_;
  assign po43 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n384_ | new_n416_ | new_n448_ | new_n480_;
  assign po44 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n385_ | new_n417_ | new_n449_ | new_n481_;
  assign po45 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n386_ | new_n418_ | new_n450_ | new_n482_;
  assign po46 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n387_ | new_n419_ | new_n451_ | new_n483_;
  assign po47 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n356_ | new_n388_ | new_n420_ | new_n452_;
  assign po48 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n357_ | new_n389_ | new_n421_ | new_n453_;
  assign po49 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n358_ | new_n390_ | new_n422_ | new_n454_;
  assign po50 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n359_ | new_n391_ | new_n423_ | new_n455_;
  assign po51 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n360_ | new_n392_ | new_n424_ | new_n456_;
  assign po52 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n361_ | new_n393_ | new_n425_ | new_n457_;
  assign po53 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n362_ | new_n394_ | new_n426_ | new_n458_;
  assign po54 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n363_ | new_n395_ | new_n427_ | new_n459_;
  assign po55 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n364_ | new_n396_ | new_n428_ | new_n460_;
  assign po56 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n365_ | new_n397_ | new_n429_ | new_n461_;
  assign po57 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n366_ | new_n398_ | new_n430_ | new_n462_;
  assign po58 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n367_ | new_n399_ | new_n431_ | new_n463_;
  assign po59 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n368_ | new_n400_ | new_n432_ | new_n464_;
  assign po60 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n369_ | new_n401_ | new_n433_ | new_n465_;
  assign po61 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n370_ | new_n402_ | new_n434_ | new_n466_;
  assign po62 = new_n498_ | new_n500_ | new_n492_ | new_n495_ | new_n371_ | new_n403_ | new_n435_ | new_n467_;
  assign new_n356_ = new_n172_ & new_n501_ & pi67 & new_n502_;
  assign new_n357_ = new_n172_ & new_n501_ & pi68 & new_n502_;
  assign new_n358_ = new_n172_ & new_n501_ & pi69 & new_n502_;
  assign new_n359_ = new_n172_ & new_n501_ & pi70 & new_n502_;
  assign new_n360_ = new_n172_ & new_n501_ & pi71 & new_n502_;
  assign new_n361_ = new_n172_ & new_n501_ & pi72 & new_n502_;
  assign new_n362_ = new_n172_ & new_n501_ & pi73 & new_n502_;
  assign new_n363_ = new_n172_ & new_n501_ & pi74 & new_n502_;
  assign new_n364_ = new_n172_ & new_n501_ & pi75 & new_n502_;
  assign new_n365_ = new_n172_ & new_n501_ & pi76 & new_n502_;
  assign new_n366_ = new_n172_ & new_n501_ & pi77 & new_n502_;
  assign new_n367_ = new_n172_ & new_n501_ & pi78 & new_n502_;
  assign new_n368_ = new_n172_ & new_n501_ & pi79 & new_n502_;
  assign new_n369_ = new_n172_ & new_n501_ & pi80 & new_n502_;
  assign new_n370_ = new_n172_ & new_n501_ & pi81 & new_n502_;
  assign new_n371_ = new_n172_ & new_n501_ & pi82 & new_n502_;
  assign new_n372_ = new_n172_ & new_n501_ & pi83 & new_n502_;
  assign new_n373_ = new_n172_ & new_n501_ & pi84 & new_n502_;
  assign new_n374_ = new_n172_ & new_n501_ & pi85 & new_n502_;
  assign new_n375_ = new_n172_ & new_n501_ & pi86 & new_n502_;
  assign new_n376_ = new_n172_ & new_n501_ & pi41 & new_n502_;
  assign new_n377_ = new_n172_ & new_n501_ & pi42 & new_n502_;
  assign new_n378_ = new_n172_ & new_n501_ & pi43 & new_n502_;
  assign new_n379_ = new_n172_ & new_n501_ & pi44 & new_n502_;
  assign new_n380_ = new_n172_ & new_n501_ & pi45 & new_n502_;
  assign new_n381_ = new_n172_ & new_n501_ & pi46 & new_n502_;
  assign new_n382_ = new_n172_ & new_n501_ & pi47 & new_n502_;
  assign new_n383_ = new_n172_ & new_n501_ & pi48 & new_n502_;
  assign new_n384_ = new_n172_ & new_n501_ & pi49 & new_n502_;
  assign new_n385_ = new_n172_ & new_n501_ & pi50 & new_n502_;
  assign new_n386_ = new_n172_ & new_n501_ & pi51 & new_n502_;
  assign new_n387_ = new_n172_ & new_n501_ & pi87 & new_n502_;
  assign new_n388_ = new_n172_ & new_n503_ & pi75 & new_n174_;
  assign new_n389_ = new_n172_ & new_n503_ & pi76 & new_n174_;
  assign new_n390_ = new_n172_ & new_n503_ & pi77 & new_n174_;
  assign new_n391_ = new_n172_ & new_n503_ & pi78 & new_n174_;
  assign new_n392_ = new_n172_ & new_n503_ & pi79 & new_n174_;
  assign new_n393_ = new_n172_ & new_n503_ & pi80 & new_n174_;
  assign new_n394_ = new_n172_ & new_n503_ & pi81 & new_n174_;
  assign new_n395_ = new_n172_ & new_n503_ & pi82 & new_n174_;
  assign new_n396_ = new_n172_ & new_n503_ & pi83 & new_n174_;
  assign new_n397_ = new_n172_ & new_n503_ & pi84 & new_n174_;
  assign new_n398_ = new_n172_ & new_n503_ & pi85 & new_n174_;
  assign new_n399_ = new_n172_ & new_n503_ & pi86 & new_n174_;
  assign new_n400_ = new_n172_ & new_n503_ & pi41 & new_n174_;
  assign new_n401_ = new_n172_ & new_n503_ & pi42 & new_n174_;
  assign new_n402_ = new_n172_ & new_n503_ & pi43 & new_n174_;
  assign new_n403_ = new_n172_ & new_n503_ & pi44 & new_n174_;
  assign new_n404_ = new_n172_ & new_n503_ & pi45 & new_n174_;
  assign new_n405_ = new_n172_ & new_n503_ & pi46 & new_n174_;
  assign new_n406_ = new_n172_ & new_n503_ & pi47 & new_n174_;
  assign new_n407_ = new_n172_ & new_n503_ & pi48 & new_n174_;
  assign new_n408_ = new_n172_ & new_n503_ & pi49 & new_n174_;
  assign new_n409_ = new_n172_ & new_n503_ & pi50 & new_n174_;
  assign new_n410_ = new_n172_ & new_n503_ & pi51 & new_n174_;
  assign new_n411_ = new_n172_ & new_n503_ & pi87 & new_n174_;
  assign new_n412_ = new_n172_ & new_n503_ & pi09 & new_n174_;
  assign new_n413_ = new_n172_ & new_n503_ & pi10 & new_n174_;
  assign new_n414_ = new_n172_ & new_n503_ & pi11 & new_n174_;
  assign new_n415_ = new_n172_ & new_n503_ & pi12 & new_n174_;
  assign new_n416_ = new_n172_ & new_n503_ & pi13 & new_n174_;
  assign new_n417_ = new_n172_ & new_n503_ & pi14 & new_n174_;
  assign new_n418_ = new_n172_ & new_n503_ & pi15 & new_n174_;
  assign new_n419_ = new_n172_ & new_n503_ & pi16 & new_n174_;
  assign new_n420_ = new_n172_ & new_n173_ & pi78 & new_n504_;
  assign new_n421_ = new_n172_ & new_n173_ & pi79 & new_n504_;
  assign new_n422_ = new_n172_ & new_n173_ & pi80 & new_n504_;
  assign new_n423_ = new_n172_ & new_n173_ & pi81 & new_n504_;
  assign new_n424_ = new_n172_ & new_n173_ & pi82 & new_n504_;
  assign new_n425_ = new_n172_ & new_n173_ & pi83 & new_n504_;
  assign new_n426_ = new_n172_ & new_n173_ & pi84 & new_n504_;
  assign new_n427_ = new_n172_ & new_n173_ & pi85 & new_n504_;
  assign new_n428_ = new_n172_ & new_n173_ & pi86 & new_n504_;
  assign new_n429_ = new_n172_ & new_n173_ & pi41 & new_n504_;
  assign new_n430_ = new_n172_ & new_n173_ & pi42 & new_n504_;
  assign new_n431_ = new_n172_ & new_n173_ & pi43 & new_n504_;
  assign new_n432_ = new_n172_ & new_n173_ & pi44 & new_n504_;
  assign new_n433_ = new_n172_ & new_n173_ & pi45 & new_n504_;
  assign new_n434_ = new_n172_ & new_n173_ & pi46 & new_n504_;
  assign new_n435_ = new_n172_ & new_n173_ & pi47 & new_n504_;
  assign new_n436_ = new_n172_ & new_n173_ & pi48 & new_n504_;
  assign new_n437_ = new_n172_ & new_n173_ & pi49 & new_n504_;
  assign new_n438_ = new_n172_ & new_n173_ & pi50 & new_n504_;
  assign new_n439_ = new_n172_ & new_n173_ & pi51 & new_n504_;
  assign new_n440_ = new_n172_ & new_n173_ & pi87 & new_n504_;
  assign new_n441_ = new_n172_ & new_n173_ & pi09 & new_n504_;
  assign new_n442_ = new_n172_ & new_n173_ & pi10 & new_n504_;
  assign new_n443_ = new_n172_ & new_n173_ & pi11 & new_n504_;
  assign new_n444_ = new_n172_ & new_n173_ & pi12 & new_n504_;
  assign new_n445_ = new_n172_ & new_n173_ & pi13 & new_n504_;
  assign new_n446_ = new_n172_ & new_n173_ & pi14 & new_n504_;
  assign new_n447_ = new_n172_ & new_n173_ & pi15 & new_n504_;
  assign new_n448_ = new_n172_ & new_n173_ & pi16 & new_n504_;
  assign new_n449_ = new_n172_ & new_n173_ & pi17 & new_n504_;
  assign new_n450_ = new_n172_ & new_n173_ & pi18 & new_n504_;
  assign new_n451_ = new_n172_ & new_n173_ & pi19 & new_n504_;
  assign new_n452_ = new_n172_ & new_n173_ & pi82 & new_n174_;
  assign new_n453_ = new_n172_ & new_n173_ & pi83 & new_n174_;
  assign new_n454_ = new_n172_ & new_n173_ & pi84 & new_n174_;
  assign new_n455_ = new_n172_ & new_n173_ & pi85 & new_n174_;
  assign new_n456_ = new_n172_ & new_n173_ & pi86 & new_n174_;
  assign new_n457_ = new_n172_ & new_n173_ & pi41 & new_n174_;
  assign new_n458_ = new_n172_ & new_n173_ & pi42 & new_n174_;
  assign new_n459_ = new_n172_ & new_n173_ & pi43 & new_n174_;
  assign new_n460_ = new_n172_ & new_n173_ & pi44 & new_n174_;
  assign new_n461_ = new_n172_ & new_n173_ & pi45 & new_n174_;
  assign new_n462_ = new_n172_ & new_n173_ & pi46 & new_n174_;
  assign new_n463_ = new_n172_ & new_n173_ & pi47 & new_n174_;
  assign new_n464_ = new_n172_ & new_n173_ & pi48 & new_n174_;
  assign new_n465_ = new_n172_ & new_n173_ & pi49 & new_n174_;
  assign new_n466_ = new_n172_ & new_n173_ & pi50 & new_n174_;
  assign new_n467_ = new_n172_ & new_n173_ & pi51 & new_n174_;
  assign new_n468_ = new_n172_ & new_n173_ & pi87 & new_n174_;
  assign new_n469_ = new_n172_ & new_n173_ & pi09 & new_n174_;
  assign new_n470_ = new_n172_ & new_n173_ & pi10 & new_n174_;
  assign new_n471_ = new_n172_ & new_n173_ & pi11 & new_n174_;
  assign new_n472_ = new_n172_ & new_n173_ & pi12 & new_n174_;
  assign new_n473_ = new_n172_ & new_n173_ & pi13 & new_n174_;
  assign new_n474_ = new_n172_ & new_n173_ & pi14 & new_n174_;
  assign new_n475_ = new_n172_ & new_n173_ & pi15 & new_n174_;
  assign new_n476_ = new_n172_ & new_n173_ & pi16 & new_n174_;
  assign new_n477_ = new_n172_ & new_n173_ & pi17 & new_n174_;
  assign new_n478_ = new_n172_ & new_n173_ & pi18 & new_n174_;
  assign new_n479_ = new_n172_ & new_n173_ & pi19 & new_n174_;
  assign new_n480_ = new_n172_ & new_n173_ & pi20 & new_n174_;
  assign new_n481_ = new_n172_ & new_n173_ & pi21 & new_n174_;
  assign new_n482_ = new_n172_ & new_n173_ & pi22 & new_n174_;
  assign new_n483_ = new_n172_ & new_n173_ & pi23 & new_n174_;
  assign new_n484_ = ~new_n173_;
  assign new_n485_ = ~new_n174_;
  assign new_n486_ = ~new_n173_;
  assign new_n487_ = new_n174_ & new_n172_ & new_n486_;
  assign new_n488_ = ~new_n174_;
  assign new_n489_ = ~new_n172_;
  assign new_n490_ = ~new_n173_;
  assign new_n491_ = ~new_n174_;
  assign new_n492_ = new_n491_ & new_n489_ & new_n490_;
  assign new_n493_ = ~new_n172_;
  assign new_n494_ = ~new_n173_;
  assign new_n495_ = new_n174_ & new_n493_ & new_n494_;
  assign new_n496_ = ~new_n172_;
  assign new_n497_ = ~new_n174_;
  assign new_n498_ = new_n497_ & new_n496_ & new_n173_;
  assign new_n499_ = ~new_n172_;
  assign new_n500_ = new_n174_ & new_n499_ & new_n173_;
  assign new_n501_ = ~new_n173_;
  assign new_n502_ = ~new_n174_;
  assign new_n503_ = ~new_n173_;
  assign new_n504_ = ~new_n174_;
endmodule


