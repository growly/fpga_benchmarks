// Benchmark "C880.iscas" written by ABC on Thu Mar 19 13:02:36 2020

module C880_iscas  ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47,
    pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45,
    pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57,
    pi58, pi59;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25;
  wire new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n161_, new_n162_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_,
    new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n183_,
    new_n184_, new_n186_, new_n187_, new_n190_, new_n192_, new_n193_,
    new_n194_, new_n196_, new_n197_, new_n198_, new_n199_, new_n201_,
    new_n202_, new_n204_, new_n205_, new_n207_, new_n208_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_,
    new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_,
    new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_,
    new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_,
    new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_,
    new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_,
    new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_,
    new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_,
    new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_,
    new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_,
    new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_,
    new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n375_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n452_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_,
    new_n459_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_;
  assign new_n87_ = ~pi59;
  assign new_n88_ = pi54 & pi58;
  assign new_n89_ = pi54 & pi56;
  assign new_n90_ = pi54 & pi55;
  assign new_n91_ = pi46 | pi47;
  assign new_n92_ = ~pi46 | ~pi47;
  assign new_n93_ = pi44 | pi45;
  assign new_n94_ = ~pi44 | ~pi45;
  assign new_n95_ = pi42 | pi43;
  assign new_n96_ = ~pi42 | ~pi43;
  assign new_n97_ = pi40 | pi41;
  assign new_n98_ = ~pi40 | ~pi41;
  assign new_n99_ = pi37 & pi33;
  assign new_n100_ = pi49 & pi29;
  assign new_n101_ = pi29 | pi30;
  assign new_n102_ = ~pi29 | ~pi30;
  assign new_n103_ = pi49 & pi28;
  assign new_n104_ = pi49 & pi27;
  assign new_n105_ = pi27 | pi28;
  assign new_n106_ = ~pi27 | ~pi28;
  assign new_n107_ = pi49 & pi26;
  assign new_n108_ = pi49 & pi25;
  assign new_n109_ = pi25 | pi26;
  assign new_n110_ = ~pi25 | ~pi26;
  assign new_n111_ = pi49 & pi24;
  assign new_n112_ = pi49 & pi23;
  assign new_n113_ = pi23 | pi24;
  assign new_n114_ = ~pi23 | ~pi24;
  assign new_n115_ = pi19 | pi20;
  assign new_n116_ = pi17 & pi18;
  assign new_n117_ = ~pi10 | ~pi39;
  assign new_n118_ = pi16 & pi10 & pi15;
  assign new_n119_ = ~pi14 | ~pi10 | ~pi11;
  assign new_n120_ = pi08 & pi33;
  assign new_n121_ = pi07 & pi10 & pi15;
  assign new_n122_ = ~pi12 | ~pi11 | ~pi10 | ~pi07;
  assign new_n123_ = pi07 & pi10 & pi06;
  assign new_n124_ = pi16 & pi10 & pi06;
  assign new_n125_ = pi07 & pi05 & pi06;
  assign new_n126_ = pi16 & pi05 & pi06;
  assign new_n127_ = pi07 & pi05 & pi15;
  assign new_n128_ = pi16 & pi05 & pi15;
  assign new_n129_ = ~pi05 | ~pi11;
  assign new_n130_ = pi07 & pi05 & pi06;
  assign new_n131_ = pi03 & pi07;
  assign new_n132_ = ~pi03 & ~pi07;
  assign new_n133_ = pi03 & pi33;
  assign new_n134_ = pi01 & pi33;
  assign new_n135_ = ~pi09 | ~pi02 | ~pi00 | ~pi01;
  assign new_n136_ = ~pi03 | ~pi08 | ~pi00 | ~pi01;
  assign new_n137_ = pi08 & pi00 & pi04;
  assign new_n138_ = ~pi03 | ~pi02 | ~pi00 | ~pi04;
  assign new_n139_ = ~pi03 | ~pi02 | ~pi00 | ~pi01;
  assign new_n140_ = ~new_n87_;
  assign new_n141_ = ~new_n92_ | ~new_n91_;
  assign new_n142_ = ~new_n94_ | ~new_n93_;
  assign new_n143_ = ~new_n96_ | ~new_n95_;
  assign new_n144_ = ~new_n98_ | ~new_n97_;
  assign new_n145_ = ~new_n102_ | ~new_n101_;
  assign new_n146_ = ~new_n106_ | ~new_n105_;
  assign new_n147_ = ~new_n110_ | ~new_n109_;
  assign new_n148_ = ~new_n114_ | ~new_n113_;
  assign new_n149_ = pi22 & new_n115_;
  assign new_n150_ = ~pi21 | ~new_n115_;
  assign po03 = new_n116_;
  assign new_n152_ = ~new_n118_;
  assign new_n153_ = new_n135_ | new_n119_;
  assign new_n154_ = ~new_n121_;
  assign new_n155_ = ~new_n135_ & ~new_n122_;
  assign new_n156_ = ~new_n123_;
  assign new_n157_ = ~new_n124_;
  assign po02 = new_n125_;
  assign po01 = new_n126_;
  assign po00 = new_n127_;
  assign new_n161_ = new_n135_ | new_n129_;
  assign new_n162_ = ~new_n130_;
  assign new_n163_ = new_n138_ | new_n130_;
  assign new_n164_ = ~new_n132_ & ~new_n131_;
  assign new_n165_ = ~new_n136_;
  assign new_n166_ = ~new_n137_;
  assign new_n167_ = ~new_n137_;
  assign new_n168_ = ~new_n139_;
  assign new_n169_ = pi49 & new_n140_;
  assign new_n170_ = ~new_n141_;
  assign new_n171_ = new_n142_ & new_n141_;
  assign new_n172_ = ~new_n142_;
  assign new_n173_ = ~new_n143_;
  assign new_n174_ = new_n144_ & new_n143_;
  assign new_n175_ = ~new_n144_;
  assign new_n176_ = ~new_n145_;
  assign new_n177_ = new_n146_ & new_n145_;
  assign new_n178_ = ~new_n146_;
  assign new_n179_ = ~new_n147_;
  assign new_n180_ = new_n148_ & new_n147_;
  assign new_n181_ = ~new_n148_;
  assign po09 = new_n149_;
  assign new_n183_ = ~new_n150_;
  assign new_n184_ = new_n155_ & pi13;
  assign po06 = new_n152_;
  assign new_n186_ = ~new_n153_;
  assign new_n187_ = ~new_n165_ | ~new_n154_;
  assign po08 = new_n156_;
  assign po07 = new_n157_;
  assign new_n190_ = ~new_n161_;
  assign po05 = new_n163_;
  assign new_n192_ = ~new_n166_;
  assign new_n193_ = ~new_n167_;
  assign new_n194_ = new_n138_ | new_n162_;
  assign po04 = new_n168_;
  assign new_n196_ = new_n172_ & new_n170_;
  assign new_n197_ = new_n175_ & new_n173_;
  assign new_n198_ = new_n178_ & new_n176_;
  assign new_n199_ = new_n181_ & new_n179_;
  assign po14 = new_n183_;
  assign new_n201_ = ~new_n184_;
  assign new_n202_ = ~new_n192_ | ~pi39 | ~new_n164_ | ~pi10;
  assign po13 = new_n186_;
  assign new_n204_ = ~pi09 | ~new_n192_ | ~new_n128_;
  assign new_n205_ = pi09 & new_n117_ & new_n192_;
  assign po12 = new_n190_;
  assign new_n207_ = ~pi03 | ~new_n192_ | ~new_n117_;
  assign new_n208_ = new_n128_ & new_n192_ & pi03;
  assign po11 = new_n193_;
  assign po10 = new_n194_;
  assign new_n211_ = new_n140_ | new_n204_;
  assign new_n212_ = new_n140_ | new_n204_;
  assign new_n213_ = new_n140_ | new_n204_;
  assign new_n214_ = new_n140_ | new_n204_;
  assign new_n215_ = new_n87_ & new_n208_;
  assign new_n216_ = new_n87_ & new_n208_;
  assign new_n217_ = new_n87_ & new_n208_;
  assign new_n218_ = new_n87_ & new_n208_;
  assign new_n219_ = ~new_n171_ & ~new_n196_;
  assign new_n220_ = ~new_n174_ & ~new_n197_;
  assign new_n221_ = pi38 & new_n205_;
  assign new_n222_ = pi36 & new_n205_;
  assign new_n223_ = pi35 & new_n205_;
  assign new_n224_ = pi34 & new_n205_;
  assign new_n225_ = ~new_n177_ & ~new_n198_;
  assign new_n226_ = ~new_n180_ & ~new_n199_;
  assign new_n227_ = ~new_n201_;
  assign new_n228_ = ~new_n202_ | ~new_n187_;
  assign new_n229_ = ~new_n207_ | ~pi00;
  assign new_n230_ = ~new_n224_ & ~new_n215_;
  assign new_n231_ = ~new_n223_ & ~new_n216_;
  assign new_n232_ = ~new_n222_ & ~new_n217_;
  assign new_n233_ = ~new_n221_ & ~new_n218_;
  assign new_n234_ = new_n219_ | pi48;
  assign new_n235_ = ~new_n219_ | ~pi48;
  assign new_n236_ = ~new_n227_ | ~pi47;
  assign new_n237_ = ~new_n227_ | ~pi46;
  assign new_n238_ = ~new_n227_ | ~pi45;
  assign new_n239_ = new_n227_ & pi44;
  assign new_n240_ = new_n227_ & pi43;
  assign new_n241_ = new_n227_ & pi42;
  assign new_n242_ = new_n227_ & pi41;
  assign new_n243_ = new_n227_ & pi40;
  assign new_n244_ = pi38 & new_n229_;
  assign new_n245_ = pi36 & new_n229_;
  assign new_n246_ = pi35 & new_n229_;
  assign new_n247_ = pi34 & new_n229_;
  assign new_n248_ = new_n225_ | pi32;
  assign new_n249_ = ~new_n225_ | ~pi32;
  assign new_n250_ = pi31 | new_n220_;
  assign new_n251_ = ~pi31 | ~new_n220_;
  assign new_n252_ = pi31 | new_n226_;
  assign new_n253_ = ~pi31 | ~new_n226_;
  assign new_n254_ = pi30 & new_n228_;
  assign new_n255_ = pi29 & new_n228_;
  assign new_n256_ = pi28 & new_n228_;
  assign new_n257_ = pi27 & new_n228_;
  assign new_n258_ = pi26 & new_n228_;
  assign new_n259_ = pi25 & new_n228_;
  assign new_n260_ = pi24 & new_n228_;
  assign new_n261_ = pi23 & new_n228_;
  assign new_n262_ = ~new_n235_ | ~new_n234_;
  assign new_n263_ = ~new_n244_ & ~new_n254_;
  assign new_n264_ = ~new_n245_ & ~new_n255_;
  assign new_n265_ = ~new_n246_ & ~new_n256_;
  assign new_n266_ = ~new_n247_ & ~new_n257_;
  assign new_n267_ = ~new_n99_ & ~new_n258_;
  assign new_n268_ = ~new_n249_ | ~new_n248_;
  assign new_n269_ = ~new_n251_ | ~new_n250_;
  assign new_n270_ = ~new_n253_ | ~new_n252_;
  assign new_n271_ = ~new_n120_ & ~new_n260_;
  assign new_n272_ = ~new_n133_ & ~new_n259_;
  assign new_n273_ = ~new_n134_ & ~new_n261_;
  assign new_n274_ = ~new_n211_ | ~new_n266_;
  assign new_n275_ = ~new_n212_ | ~new_n265_;
  assign new_n276_ = ~new_n213_ | ~new_n264_;
  assign new_n277_ = ~new_n214_ | ~new_n263_;
  assign new_n278_ = ~new_n273_ | ~new_n230_;
  assign new_n279_ = ~new_n271_ | ~new_n231_;
  assign new_n280_ = ~new_n272_ | ~new_n232_;
  assign new_n281_ = ~new_n267_ | ~new_n233_;
  assign new_n282_ = ~new_n262_;
  assign new_n283_ = new_n269_ & new_n262_;
  assign new_n284_ = ~new_n268_;
  assign new_n285_ = new_n270_ & new_n268_;
  assign new_n286_ = ~new_n269_;
  assign new_n287_ = ~new_n270_;
  assign new_n288_ = pi53 & new_n277_;
  assign new_n289_ = pi53 & new_n276_;
  assign new_n290_ = pi53 & new_n275_;
  assign new_n291_ = pi53 & new_n274_;
  assign new_n292_ = pi53 & new_n281_;
  assign new_n293_ = pi53 & new_n280_;
  assign new_n294_ = pi53 & new_n279_;
  assign new_n295_ = pi53 & new_n278_;
  assign new_n296_ = new_n286_ & new_n282_;
  assign new_n297_ = new_n277_ | pi47;
  assign new_n298_ = ~new_n277_ | ~pi47;
  assign new_n299_ = new_n276_ | pi46;
  assign new_n300_ = ~new_n276_ | ~pi46;
  assign new_n301_ = new_n275_ | pi45;
  assign new_n302_ = ~new_n275_ | ~pi45;
  assign new_n303_ = new_n274_ | pi44;
  assign new_n304_ = ~new_n274_ | ~pi44;
  assign new_n305_ = new_n281_ | pi43;
  assign new_n306_ = ~new_n281_ | ~pi43;
  assign new_n307_ = new_n280_ | pi42;
  assign new_n308_ = ~new_n280_ | ~pi42;
  assign new_n309_ = new_n279_ | pi41;
  assign new_n310_ = ~new_n279_ | ~pi41;
  assign new_n311_ = new_n278_ | pi40;
  assign new_n312_ = ~new_n278_ | ~pi40;
  assign new_n313_ = new_n287_ & new_n284_;
  assign new_n314_ = ~pi57 | ~new_n297_ | ~new_n301_ | ~new_n299_;
  assign new_n315_ = ~pi57 | ~new_n299_ | ~new_n297_;
  assign new_n316_ = ~new_n297_ | ~pi57;
  assign new_n317_ = ~new_n88_ & ~new_n288_;
  assign new_n318_ = ~new_n89_ & ~new_n289_;
  assign new_n319_ = ~new_n90_ & ~new_n290_;
  assign new_n320_ = ~new_n283_ & ~new_n296_;
  assign new_n321_ = new_n297_ & new_n298_;
  assign new_n322_ = ~new_n298_;
  assign new_n323_ = new_n299_ & new_n300_;
  assign new_n324_ = ~new_n300_;
  assign new_n325_ = new_n301_ & new_n302_;
  assign new_n326_ = ~new_n302_;
  assign new_n327_ = new_n303_ & new_n304_;
  assign new_n328_ = ~new_n304_;
  assign new_n329_ = ~new_n291_ & ~new_n239_;
  assign new_n330_ = new_n305_ & new_n306_;
  assign new_n331_ = ~new_n306_;
  assign new_n332_ = ~new_n292_ & ~new_n240_;
  assign new_n333_ = new_n307_ & new_n308_;
  assign new_n334_ = ~new_n308_;
  assign new_n335_ = ~new_n293_ & ~new_n241_;
  assign new_n336_ = new_n309_ & new_n310_;
  assign new_n337_ = ~new_n310_;
  assign new_n338_ = ~new_n294_ & ~new_n242_;
  assign new_n339_ = new_n311_ & new_n312_;
  assign new_n340_ = ~new_n312_;
  assign new_n341_ = ~new_n295_ & ~new_n243_;
  assign new_n342_ = ~new_n285_ & ~new_n313_;
  assign new_n343_ = new_n321_ & pi57;
  assign new_n344_ = ~new_n321_ & ~pi57;
  assign new_n345_ = pi52 & new_n322_;
  assign new_n346_ = pi52 & new_n324_;
  assign new_n347_ = pi52 & new_n326_;
  assign new_n348_ = pi52 & new_n328_;
  assign new_n349_ = pi52 & new_n331_;
  assign new_n350_ = pi52 & new_n334_;
  assign new_n351_ = pi52 & new_n337_;
  assign new_n352_ = pi52 & new_n340_;
  assign new_n353_ = pi51 & new_n321_;
  assign new_n354_ = pi51 & new_n323_;
  assign new_n355_ = pi51 & new_n325_;
  assign new_n356_ = pi51 & new_n327_;
  assign new_n357_ = pi51 & new_n330_;
  assign new_n358_ = pi51 & new_n333_;
  assign new_n359_ = pi51 & new_n336_;
  assign new_n360_ = pi51 & new_n339_;
  assign po16 = new_n320_;
  assign new_n362_ = ~new_n322_;
  assign new_n363_ = ~new_n299_ | ~new_n322_;
  assign new_n364_ = ~new_n322_ | ~new_n301_ | ~new_n299_;
  assign new_n365_ = ~new_n324_;
  assign new_n366_ = ~new_n301_ | ~new_n324_;
  assign new_n367_ = ~new_n326_;
  assign new_n368_ = ~new_n328_;
  assign new_n369_ = ~new_n331_;
  assign new_n370_ = ~new_n307_ | ~new_n331_;
  assign new_n371_ = ~new_n331_ | ~new_n309_ | ~new_n307_;
  assign new_n372_ = ~new_n334_;
  assign new_n373_ = ~new_n309_ | ~new_n334_;
  assign new_n374_ = ~new_n337_;
  assign new_n375_ = ~new_n340_;
  assign po15 = new_n342_;
  assign new_n377_ = ~new_n344_ & ~new_n343_;
  assign new_n378_ = ~new_n314_ | ~new_n364_ | ~new_n367_ | ~new_n366_;
  assign new_n379_ = ~new_n315_ | ~new_n365_ | ~new_n363_;
  assign new_n380_ = ~new_n362_ | ~new_n316_;
  assign new_n381_ = ~new_n353_ & ~new_n345_;
  assign new_n382_ = ~new_n354_ & ~new_n346_;
  assign new_n383_ = ~new_n355_ & ~new_n347_;
  assign new_n384_ = ~new_n356_ & ~new_n348_;
  assign new_n385_ = ~new_n357_ & ~new_n349_;
  assign new_n386_ = ~new_n358_ & ~new_n350_;
  assign new_n387_ = ~new_n359_ & ~new_n351_;
  assign new_n388_ = ~new_n360_ & ~new_n352_;
  assign new_n389_ = pi50 & new_n377_;
  assign new_n390_ = ~new_n323_ & ~new_n380_;
  assign new_n391_ = new_n323_ & new_n380_;
  assign new_n392_ = ~new_n325_ & ~new_n379_;
  assign new_n393_ = new_n325_ & new_n379_;
  assign new_n394_ = ~new_n327_ & ~new_n378_;
  assign new_n395_ = new_n327_ & new_n378_;
  assign new_n396_ = ~new_n303_ | ~new_n378_;
  assign new_n397_ = ~new_n390_ & ~new_n391_;
  assign new_n398_ = ~new_n392_ & ~new_n393_;
  assign new_n399_ = ~new_n394_ & ~new_n395_;
  assign new_n400_ = ~new_n396_ | ~new_n368_;
  assign new_n401_ = ~new_n100_ & ~new_n389_;
  assign new_n402_ = pi50 & new_n397_;
  assign new_n403_ = pi50 & new_n398_;
  assign new_n404_ = pi50 & new_n399_;
  assign new_n405_ = ~new_n236_ | ~new_n317_ | ~new_n401_ | ~new_n381_;
  assign new_n406_ = ~new_n330_ & ~new_n400_;
  assign new_n407_ = new_n330_ & new_n400_;
  assign new_n408_ = ~new_n305_ | ~new_n400_;
  assign new_n409_ = ~new_n400_ | ~new_n307_ | ~new_n305_;
  assign new_n410_ = ~new_n400_ | ~new_n305_ | ~new_n309_ | ~new_n307_;
  assign new_n411_ = ~new_n405_;
  assign new_n412_ = ~new_n406_ & ~new_n407_;
  assign new_n413_ = ~new_n369_ | ~new_n408_;
  assign new_n414_ = ~new_n409_ | ~new_n372_ | ~new_n370_;
  assign new_n415_ = ~new_n410_ | ~new_n371_ | ~new_n374_ | ~new_n373_;
  assign new_n416_ = ~new_n103_ & ~new_n402_;
  assign new_n417_ = ~new_n104_ & ~new_n403_;
  assign new_n418_ = ~new_n107_ & ~new_n404_;
  assign new_n419_ = pi50 & new_n412_;
  assign new_n420_ = ~new_n411_;
  assign new_n421_ = ~new_n237_ | ~new_n318_ | ~new_n416_ | ~new_n382_;
  assign new_n422_ = ~new_n238_ | ~new_n319_ | ~new_n417_ | ~new_n383_;
  assign new_n423_ = ~new_n329_ | ~new_n418_ | ~new_n384_;
  assign new_n424_ = ~new_n333_ & ~new_n413_;
  assign new_n425_ = new_n333_ & new_n413_;
  assign new_n426_ = ~new_n336_ & ~new_n414_;
  assign new_n427_ = new_n336_ & new_n414_;
  assign new_n428_ = ~new_n339_ & ~new_n415_;
  assign new_n429_ = new_n339_ & new_n415_;
  assign new_n430_ = ~new_n415_ | ~new_n311_;
  assign po17 = new_n420_;
  assign new_n432_ = ~new_n421_;
  assign new_n433_ = ~new_n422_;
  assign new_n434_ = ~new_n423_;
  assign new_n435_ = ~new_n424_ & ~new_n425_;
  assign new_n436_ = ~new_n426_ & ~new_n427_;
  assign new_n437_ = ~new_n428_ & ~new_n429_;
  assign new_n438_ = new_n375_ & new_n430_;
  assign new_n439_ = ~new_n108_ & ~new_n419_;
  assign new_n440_ = pi50 & new_n435_;
  assign new_n441_ = pi50 & new_n436_;
  assign new_n442_ = pi50 & new_n437_;
  assign new_n443_ = ~new_n432_;
  assign new_n444_ = ~new_n433_;
  assign new_n445_ = ~new_n434_;
  assign new_n446_ = ~new_n332_ | ~new_n439_ | ~new_n385_;
  assign new_n447_ = ~new_n438_;
  assign new_n448_ = ~new_n169_ & ~new_n442_;
  assign po20 = new_n443_;
  assign po19 = new_n444_;
  assign po18 = new_n445_;
  assign new_n452_ = ~new_n446_;
  assign po21 = new_n447_;
  assign new_n454_ = ~new_n111_ & ~new_n440_;
  assign new_n455_ = ~new_n112_ & ~new_n441_;
  assign new_n456_ = ~new_n452_;
  assign new_n457_ = ~new_n335_ | ~new_n454_ | ~new_n386_;
  assign new_n458_ = ~new_n338_ | ~new_n455_ | ~new_n387_;
  assign new_n459_ = ~new_n341_ | ~new_n448_ | ~new_n388_;
  assign po22 = new_n456_;
  assign new_n461_ = ~new_n457_;
  assign new_n462_ = ~new_n458_;
  assign new_n463_ = ~new_n459_;
  assign new_n464_ = ~new_n461_;
  assign new_n465_ = ~new_n462_;
  assign new_n466_ = ~new_n463_;
  assign po25 = new_n464_;
  assign po24 = new_n465_;
  assign po23 = new_n466_;
endmodule


