// Benchmark "frg2" written by ABC on Thu Mar 19 13:02:36 2020

module frg2 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138;
  wire new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_;
  assign po000 = ~pi057;
  assign po001 = ~new_n750_ & ((~new_n748_ & (~pi036 | ~new_n749_)) | ~pi038 | (pi036 & ~new_n749_));
  assign po002 = ~new_n753_ & ((~new_n751_ & (~pi036 | ~new_n752_)) | ~pi038 | (pi036 & ~new_n752_));
  assign po003 = ~new_n756_ & ((~new_n754_ & (~pi036 | ~new_n755_)) | ~pi038 | (pi036 & ~new_n755_));
  assign po004 = ~new_n759_ & ((~new_n757_ & (~pi036 | ~new_n758_)) | ~pi038 | (pi036 & ~new_n758_));
  assign po007 = ~new_n760_ & ((pi036 & pi037) | pi115 | (~pi036 & ~pi037));
  assign po008 = ~new_n761_ & ((pi036 & pi037) | pi116 | (~pi036 & ~pi037));
  assign po009 = ~new_n762_ & ((pi036 & pi037) | pi117 | (~pi036 & ~pi037));
  assign po010 = ~new_n763_ & ((pi036 & pi037) | pi118 | (~pi036 & ~pi037));
  assign po011 = ~new_n764_ & ((pi036 & pi037) | pi119 | (~pi036 & ~pi037));
  assign po012 = ~new_n765_ & ((pi036 & pi037) | pi120 | (~pi036 & ~pi037));
  assign po013 = ~new_n766_ & ((pi036 & pi037) | pi121 | (~pi036 & ~pi037));
  assign po014 = ~new_n767_ & ((pi036 & pi037) | pi122 | (~pi036 & ~pi037));
  assign po015 = pi115 & pi038;
  assign po016 = pi116 & pi038;
  assign po017 = pi117 & pi038;
  assign po018 = pi118 & pi038;
  assign po019 = pi119 & pi038;
  assign po020 = pi120 & pi038;
  assign po021 = pi121 & pi038;
  assign po022 = pi122 & pi038;
  assign po023 = ~pi138 & pi057;
  assign po025 = ~new_n768_;
  assign po026 = ~new_n769_;
  assign po027 = ~new_n770_;
  assign po028 = ~new_n771_;
  assign po029 = ~new_n772_;
  assign po030 = (pi064 | ~new_n775_) & (~new_n682_ | ~new_n773_ | ~new_n774_);
  assign po031 = (pi064 | ~new_n775_) & (~new_n682_ | ~new_n773_ | ~new_n774_);
  assign po032 = (pi064 | ~new_n775_) & (~new_n682_ | ~new_n773_ | ~new_n774_);
  assign po033 = (pi064 | ~new_n775_) & (~new_n682_ | ~new_n773_ | ~new_n774_);
  assign po034 = (pi064 | ~new_n775_) & (~new_n682_ | ~new_n773_ | ~new_n774_);
  assign po035 = ~new_n776_;
  assign po036 = ~new_n777_;
  assign po037 = ~new_n778_;
  assign po038 = ~new_n779_;
  assign po039 = ~new_n780_;
  assign po040 = ~new_n781_;
  assign po041 = ~new_n782_;
  assign po042 = ~new_n783_;
  assign po043 = ~new_n784_;
  assign po044 = ~new_n785_;
  assign po045 = ~pi058;
  assign po046 = ~pi059;
  assign po047 = ~pi060;
  assign po048 = ~pi061;
  assign po049 = ~pi062;
  assign po051 = ~pi056 ^ pi137;
  assign po052 = ~new_n786_ & ~pi131 & ~pi130;
  assign po053 = pi040 & ~new_n418_ & ~pi042;
  assign po054 = (pi040 & ~new_n421_ & ~new_n422_) | (~pi039 & ~new_n419_ & ~new_n420_);
  assign po055 = ~new_n427_ & (~pi057 | ~new_n426_) & (~new_n424_ | pi039 | ~new_n425_);
  assign po056 = ~new_n430_ & (~pi057 | ~new_n426_) & (~new_n424_ | pi039 | ~new_n429_);
  assign po057 = ~new_n433_ & (~pi057 | ~new_n426_) & (~new_n424_ | pi039 | ~new_n432_);
  assign po058 = ~new_n436_ & (~new_n435_ | (~pi057 & pi062));
  assign po059 = ~new_n438_ & (pi063 | (~pi039 & pi041));
  assign po060 = ~new_n442_ & (pi064 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n439_ | ~new_n440_);
  assign po061 = ~new_n447_ & (pi065 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n446_ | ~new_n440_);
  assign po062 = ~new_n450_ & (pi066 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n449_ | ~new_n440_);
  assign po063 = ~new_n453_ & (pi067 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n452_ | ~new_n440_);
  assign po064 = ~new_n456_ & (pi068 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n455_ | ~new_n440_);
  assign po065 = ~new_n459_ & (pi069 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n458_ | ~new_n440_);
  assign po066 = ~new_n462_ & (pi070 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n461_ | ~new_n440_);
  assign po067 = ~new_n465_ & (pi071 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n464_ | ~new_n440_);
  assign po068 = ~new_n468_ & (pi072 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n467_ | ~new_n440_);
  assign po069 = ~new_n471_ & (pi073 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n470_ | ~new_n440_);
  assign po070 = ~new_n474_ & (pi074 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n473_ | ~new_n440_);
  assign po071 = ~new_n477_ & (pi075 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n476_ | ~new_n440_);
  assign po072 = ~new_n480_ & (pi076 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n479_ | ~new_n440_);
  assign po073 = ~new_n483_ & (pi077 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n482_ | ~new_n440_);
  assign po074 = ~new_n486_ & (pi078 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n485_ | ~new_n440_);
  assign po075 = ~new_n489_ & (pi079 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n488_ | ~new_n440_);
  assign po076 = ~new_n492_ & (pi080 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n491_ | ~new_n440_);
  assign po077 = ~new_n495_ & (pi081 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n494_ | ~new_n440_);
  assign po078 = ~new_n498_ & (pi082 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n497_ | ~new_n440_);
  assign po079 = ~new_n501_ & (pi083 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n500_ | ~new_n440_);
  assign po080 = ~new_n504_ & (pi084 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n503_ | ~new_n440_);
  assign po081 = ~new_n507_ & (pi085 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n506_ | ~new_n440_);
  assign po082 = ~new_n510_ & (pi086 | ~pi039 | ~new_n441_) & (new_n445_ | ~new_n509_ | ~new_n440_);
  assign po083 = ~new_n512_ & ~pi042 & pi040;
  assign po084 = ~new_n517_ & ~pi042 & pi040;
  assign po085 = ~new_n521_ & ~pi042 & pi040;
  assign po086 = ~new_n525_ & ~pi042 & pi040;
  assign po087 = ~new_n529_ & ~pi042 & pi040;
  assign po088 = ~new_n533_ & ~pi042 & pi040;
  assign po089 = ~new_n537_ & ~pi042 & pi040;
  assign po090 = ~new_n541_ & ~pi042 & pi040;
  assign po091 = ~new_n545_ & ~pi042 & pi040;
  assign po092 = ~new_n554_ & ~pi042 & pi040;
  assign po093 = ~new_n557_ & ~pi042 & pi040;
  assign po094 = ~new_n560_ & ~pi042 & pi040;
  assign po095 = ~new_n563_ & ~pi042 & pi040;
  assign po096 = ~new_n566_ & ~pi042 & pi040;
  assign po097 = ~new_n569_ & ~pi042 & pi040;
  assign po098 = (pi040 & ~new_n574_ & ~new_n575_) | (~new_n572_ & ~new_n573_ & ~new_n550_);
  assign po099 = (pi040 & ~new_n579_ & ~new_n580_) | (~new_n576_ & ~new_n577_ & ~new_n578_);
  assign po100 = (pi040 & ~new_n597_ & ~new_n580_) | (~new_n576_ & ~new_n596_ & ~new_n578_);
  assign po101 = (pi040 & ~new_n599_ & ~new_n580_) | (~new_n576_ & ~new_n598_ & ~new_n578_);
  assign po102 = (pi040 & ~new_n601_ & ~new_n580_) | (~new_n576_ & ~new_n600_ & ~new_n578_);
  assign po103 = (pi040 & ~new_n603_ & ~new_n580_) | (~new_n576_ & ~new_n602_ & ~new_n578_);
  assign po104 = (pi040 & ~new_n605_ & ~new_n580_) | (~new_n576_ & ~new_n604_ & ~new_n578_);
  assign po105 = (pi040 & ~new_n607_ & ~new_n580_) | (~new_n576_ & ~new_n606_ & ~new_n578_);
  assign po106 = (pi040 & ~new_n609_ & ~new_n580_) | (~new_n576_ & ~new_n608_ & ~new_n578_);
  assign po107 = (pi040 & ~new_n611_ & ~new_n580_) | (~new_n576_ & ~new_n610_ & ~new_n578_);
  assign po108 = (pi040 & ~new_n613_ & ~new_n580_) | (~new_n576_ & ~new_n612_ & ~new_n578_);
  assign po109 = (pi040 & ~new_n615_ & ~new_n580_) | (~new_n576_ & ~new_n614_ & ~new_n578_);
  assign po110 = (pi040 & ~new_n617_ & ~new_n580_) | (~new_n576_ & ~new_n616_ & ~new_n578_);
  assign po111 = (pi040 & ~new_n619_ & ~new_n580_) | (~new_n576_ & ~new_n618_ & ~new_n578_);
  assign po112 = (pi040 & ~new_n621_ & ~new_n580_) | (~new_n576_ & ~new_n620_ & ~new_n578_);
  assign po113 = (pi040 & ~new_n623_ & ~new_n580_) | (~new_n576_ & ~new_n622_ & ~new_n578_);
  assign po114 = (pi040 & ~new_n625_ & ~new_n580_) | (~new_n576_ & ~new_n624_ & ~new_n578_);
  assign po115 = (pi040 & ~new_n627_ & ~new_n580_) | (~new_n576_ & ~new_n626_ & ~new_n578_);
  assign po116 = (pi040 & ~new_n629_ & ~new_n580_) | (~new_n576_ & ~new_n628_ & ~new_n578_);
  assign po117 = (pi040 & ~new_n631_ & ~new_n580_) | (~new_n576_ & ~new_n630_ & ~new_n578_);
  assign po118 = (pi040 & ~new_n633_ & ~new_n580_) | (~new_n576_ & ~new_n632_ & ~new_n578_);
  assign po119 = (pi040 & ~new_n635_ & ~new_n580_) | (~new_n576_ & ~new_n634_ & ~new_n578_);
  assign po120 = (pi040 & ~new_n637_ & ~new_n580_) | (~new_n576_ & ~new_n636_ & ~new_n578_);
  assign po121 = (pi040 & ~new_n641_ & ~new_n642_) | (~new_n638_ & ~new_n639_ & ~new_n640_);
  assign po122 = ~new_n653_ & (pi126 | (pi140 & ~new_n445_));
  assign po123 = ~new_n656_ | ~pi040 | (pi127 & ~new_n655_);
  assign po124 = ~new_n660_ | ~pi040 | (pi128 & ~new_n659_);
  assign po125 = ~new_n664_ & ~pi042 & pi040;
  assign po126 = ~new_n678_ | (pi040 & ~new_n676_ & ~new_n677_) | (~new_n673_ & ~new_n674_ & ~new_n675_);
  assign po127 = ~new_n687_ | (pi040 & ~new_n685_ & ~new_n686_) | (~new_n684_ & ~new_n674_ & ~new_n675_);
  assign po128 = pi040 & ((~new_n693_ & ~new_n694_) | (~pi039 & ~new_n695_));
  assign po129 = ~new_n699_ | ~pi040 | (pi133 & ~new_n698_);
  assign po130 = ~new_n704_ | ~pi040 | (pi134 & ~new_n703_);
  assign po131 = ~new_n713_ | (pi040 & ~new_n711_ & ~new_n712_) | (~new_n709_ & ~new_n710_ & ~new_n675_);
  assign po132 = ~new_n678_ | (pi040 & ~new_n720_ & ~new_n721_) | (~new_n719_ & ~new_n576_ & ~new_n675_);
  assign po133 = pi140 & ~new_n727_ & (pi137 | pi064);
  assign po134 = (pi040 & ~new_n731_ & ~new_n732_) | (~new_n729_ & ~new_n730_ & ~new_n640_);
  assign po135 = ~new_n743_ & ~pi131 & ~pi130;
  assign po136 = pi063 & ~new_n745_;
  assign po137 = ~new_n747_ & (~new_n418_ | ~new_n746_);
  assign po138 = pi139 & ~new_n576_;
  assign new_n418_ = ~new_n794_ | (~new_n793_ & ((~pi048 & pi058) | (~pi049 & pi059)));
  assign new_n419_ = ~pi040 | pi053 | pi042;
  assign new_n420_ = pi054 | ~new_n424_ | pi055;
  assign new_n421_ = pi042 | ~pi058 | pi057;
  assign new_n422_ = ~new_n423_ & new_n424_ & ~pi039;
  assign new_n423_ = pi055 & (pi054 | pi053);
  assign new_n424_ = ~new_n802_ & ~pi062 & ~pi061;
  assign new_n425_ = (~pi053 & (~pi054 | ~pi055)) | (pi054 & ~pi055);
  assign new_n426_ = pi039 | ~new_n424_ | pi055;
  assign new_n427_ = ~new_n428_ | pi042 | ~pi040;
  assign new_n428_ = pi059 | (~pi039 & ~pi055 & new_n424_);
  assign new_n429_ = (~pi054 & (~pi053 | ~pi055)) | (pi053 & ~pi055);
  assign new_n430_ = ~new_n431_ | pi042 | ~pi040;
  assign new_n431_ = pi060 | (~pi039 & ~pi055 & new_n424_);
  assign new_n432_ = (~pi054 & ~pi055) | (~pi053 & (~pi054 | ~pi055));
  assign new_n433_ = ~new_n434_ | pi042 | ~pi040;
  assign new_n434_ = pi061 | (~pi039 & ~pi055 & new_n424_);
  assign new_n435_ = ~new_n437_ | pi053 | pi039;
  assign new_n436_ = ~pi040 | pi042 | (~pi039 & ~pi055 & new_n424_);
  assign new_n437_ = new_n424_ & ~pi054;
  assign new_n438_ = ~pi040 | pi042 | (~new_n418_ & pi063);
  assign new_n439_ = pi140 & ~pi065;
  assign new_n440_ = ~new_n424_ | pi039;
  assign new_n441_ = ~pi140 | new_n445_;
  assign new_n442_ = ~new_n444_ | (~pi064 & ~new_n424_ & ~new_n443_);
  assign new_n443_ = pi140 & ~new_n445_;
  assign new_n444_ = pi040 & ~pi042 & (pi035 | pi039 | ~new_n424_);
  assign new_n445_ = ~new_n803_ & ~pi131 & ~pi130;
  assign new_n446_ = pi140 & ~pi066;
  assign new_n447_ = ~new_n448_ | (~pi065 & ~new_n424_ & ~new_n443_);
  assign new_n448_ = pi040 & ~pi042 & (pi034 | pi039 | ~new_n424_);
  assign new_n449_ = pi140 & ~pi067;
  assign new_n450_ = ~new_n451_ | (~pi066 & ~new_n424_ & ~new_n443_);
  assign new_n451_ = pi040 & ~pi042 & (pi033 | pi039 | ~new_n424_);
  assign new_n452_ = pi140 & ~pi068;
  assign new_n453_ = ~new_n454_ | (~pi067 & ~new_n424_ & ~new_n443_);
  assign new_n454_ = pi040 & ~pi042 & (pi032 | pi039 | ~new_n424_);
  assign new_n455_ = pi140 & ~pi069;
  assign new_n456_ = ~new_n457_ | (~pi068 & ~new_n424_ & ~new_n443_);
  assign new_n457_ = pi040 & ~pi042 & (pi031 | pi039 | ~new_n424_);
  assign new_n458_ = pi140 & ~pi070;
  assign new_n459_ = ~new_n460_ | (~pi069 & ~new_n424_ & ~new_n443_);
  assign new_n460_ = pi040 & ~pi042 & (pi030 | pi039 | ~new_n424_);
  assign new_n461_ = pi140 & ~pi071;
  assign new_n462_ = ~new_n463_ | (~pi070 & ~new_n424_ & ~new_n443_);
  assign new_n463_ = pi040 & ~pi042 & (pi029 | pi039 | ~new_n424_);
  assign new_n464_ = pi140 & ~pi072;
  assign new_n465_ = ~new_n466_ | (~pi071 & ~new_n424_ & ~new_n443_);
  assign new_n466_ = pi040 & ~pi042 & (pi038 | pi039 | ~new_n424_);
  assign new_n467_ = pi140 & ~pi073;
  assign new_n468_ = ~new_n469_ | (~pi072 & ~new_n424_ & ~new_n443_);
  assign new_n469_ = pi040 & ~pi042 & (pi036 | pi039 | ~new_n424_);
  assign new_n470_ = pi140 & ~pi074;
  assign new_n471_ = ~new_n472_ | (~pi073 & ~new_n424_ & ~new_n443_);
  assign new_n472_ = pi040 & ~pi042 & (pi037 | pi039 | ~new_n424_);
  assign new_n473_ = pi140 & ~pi075;
  assign new_n474_ = ~new_n475_ | (~pi074 & ~new_n424_ & ~new_n443_);
  assign new_n475_ = pi040 & ~pi042 & (pi016 | pi039 | ~new_n424_);
  assign new_n476_ = pi140 & ~pi076;
  assign new_n477_ = ~new_n478_ | (~pi075 & ~new_n424_ & ~new_n443_);
  assign new_n478_ = pi040 & ~pi042 & (pi017 | pi039 | ~new_n424_);
  assign new_n479_ = pi140 & ~pi077;
  assign new_n480_ = ~new_n481_ | (~pi076 & ~new_n424_ & ~new_n443_);
  assign new_n481_ = pi040 & ~pi042 & (pi018 | pi039 | ~new_n424_);
  assign new_n482_ = pi140 & ~pi078;
  assign new_n483_ = ~new_n484_ | (~pi077 & ~new_n424_ & ~new_n443_);
  assign new_n484_ = pi040 & ~pi042 & (pi019 | pi039 | ~new_n424_);
  assign new_n485_ = pi140 & ~pi079;
  assign new_n486_ = ~new_n487_ | (~pi078 & ~new_n424_ & ~new_n443_);
  assign new_n487_ = pi040 & ~pi042 & (pi020 | pi039 | ~new_n424_);
  assign new_n488_ = pi140 & ~pi080;
  assign new_n489_ = ~new_n490_ | (~pi079 & ~new_n424_ & ~new_n443_);
  assign new_n490_ = pi040 & ~pi042 & (pi021 | pi039 | ~new_n424_);
  assign new_n491_ = pi140 & ~pi081;
  assign new_n492_ = ~new_n493_ | (~pi080 & ~new_n424_ & ~new_n443_);
  assign new_n493_ = pi040 & ~pi042 & (pi022 | pi039 | ~new_n424_);
  assign new_n494_ = pi140 & ~pi082;
  assign new_n495_ = ~new_n496_ | (~pi081 & ~new_n424_ & ~new_n443_);
  assign new_n496_ = pi040 & ~pi042 & (pi023 | pi039 | ~new_n424_);
  assign new_n497_ = pi140 & ~pi083;
  assign new_n498_ = ~new_n499_ | (~pi082 & ~new_n424_ & ~new_n443_);
  assign new_n499_ = pi040 & ~pi042 & (pi024 | pi039 | ~new_n424_);
  assign new_n500_ = pi140 & ~pi084;
  assign new_n501_ = ~new_n502_ | (~pi083 & ~new_n424_ & ~new_n443_);
  assign new_n502_ = pi040 & ~pi042 & (pi025 | pi039 | ~new_n424_);
  assign new_n503_ = pi140 & ~pi085;
  assign new_n504_ = ~new_n505_ | (~pi084 & ~new_n424_ & ~new_n443_);
  assign new_n505_ = pi040 & ~pi042 & (pi026 | pi039 | ~new_n424_);
  assign new_n506_ = pi140 & ~pi086;
  assign new_n507_ = ~new_n508_ | (~pi085 & ~new_n424_ & ~new_n443_);
  assign new_n508_ = pi040 & ~pi042 & (pi027 | pi039 | ~new_n424_);
  assign new_n509_ = pi140 & ~pi087;
  assign new_n510_ = ~new_n511_ | (~pi086 & ~new_n424_ & ~new_n443_);
  assign new_n511_ = pi040 & ~pi042 & (pi028 | pi039 | ~new_n424_);
  assign new_n512_ = ~new_n516_ | (~pi038 & ~new_n440_ & ~new_n513_) | (~new_n445_ & ~new_n514_ & ~new_n515_);
  assign new_n513_ = (pi036 & ~pi037 & pi008) | (pi000 & (~pi036 | pi037));
  assign new_n514_ = ~pi140 | pi088;
  assign new_n515_ = ~pi038 & new_n424_ & ~pi039;
  assign new_n516_ = pi087 | (~new_n445_ & pi140) | (~pi038 & ~pi039 & new_n424_);
  assign new_n517_ = ~new_n520_ | (~pi038 & ~new_n440_ & ~new_n518_) | (~new_n445_ & ~new_n519_ & ~new_n515_);
  assign new_n518_ = (pi036 & ~pi037 & pi009) | (pi001 & (~pi036 | pi037));
  assign new_n519_ = ~pi140 | pi089;
  assign new_n520_ = pi088 | (~new_n445_ & pi140) | (~pi038 & ~pi039 & new_n424_);
  assign new_n521_ = ~new_n524_ | (~pi038 & ~new_n440_ & ~new_n522_) | (~new_n445_ & ~new_n523_ & ~new_n515_);
  assign new_n522_ = (pi036 & ~pi037 & pi010) | (pi002 & (~pi036 | pi037));
  assign new_n523_ = ~pi140 | pi090;
  assign new_n524_ = pi089 | (~new_n445_ & pi140) | (~pi038 & ~pi039 & new_n424_);
  assign new_n525_ = ~new_n528_ | (~pi038 & ~new_n440_ & ~new_n526_) | (~new_n445_ & ~new_n527_ & ~new_n515_);
  assign new_n526_ = (pi036 & ~pi037 & pi011) | (pi003 & (~pi036 | pi037));
  assign new_n527_ = ~pi140 | pi091;
  assign new_n528_ = pi090 | (~new_n445_ & pi140) | (~pi038 & ~pi039 & new_n424_);
  assign new_n529_ = ~new_n532_ | (~pi038 & ~new_n440_ & ~new_n530_) | (~new_n445_ & ~new_n531_ & ~new_n515_);
  assign new_n530_ = (pi036 & ~pi037 & pi012) | (pi004 & (~pi036 | pi037));
  assign new_n531_ = ~pi140 | pi092;
  assign new_n532_ = pi091 | (~new_n445_ & pi140) | (~pi038 & ~pi039 & new_n424_);
  assign new_n533_ = ~new_n536_ | (~pi038 & ~new_n440_ & ~new_n534_) | (~new_n445_ & ~new_n535_ & ~new_n515_);
  assign new_n534_ = (pi036 & ~pi037 & pi013) | (pi005 & (~pi036 | pi037));
  assign new_n535_ = ~pi140 | pi093;
  assign new_n536_ = pi092 | (~new_n445_ & pi140) | (~pi038 & ~pi039 & new_n424_);
  assign new_n537_ = ~new_n540_ | (~pi038 & ~new_n440_ & ~new_n538_) | (~new_n445_ & ~new_n539_ & ~new_n515_);
  assign new_n538_ = (pi036 & ~pi037 & pi014) | (pi006 & (~pi036 | pi037));
  assign new_n539_ = ~pi140 | pi094;
  assign new_n540_ = pi093 | (~new_n445_ & pi140) | (~pi038 & ~pi039 & new_n424_);
  assign new_n541_ = ~new_n544_ | (~pi038 & ~new_n440_ & ~new_n542_) | (~new_n445_ & ~new_n543_ & ~new_n515_);
  assign new_n542_ = (pi036 & ~pi037 & pi015) | (pi007 & (~pi036 | pi037));
  assign new_n543_ = ~pi140 | pi095;
  assign new_n544_ = pi094 | (~new_n445_ & pi140) | (~pi038 & ~pi039 & new_n424_);
  assign new_n545_ = ~new_n548_ & ((~pi095 & (new_n445_ | ~new_n546_)) | ~new_n547_ | (~new_n445_ & ~new_n546_));
  assign new_n546_ = pi140 & pi096;
  assign new_n547_ = ~new_n553_ | pi039 | pi038;
  assign new_n548_ = (~pi140 & pi095 & ~new_n551_) | (pi008 & ~new_n549_ & ~new_n550_);
  assign new_n549_ = pi038 | ~new_n424_ | pi039;
  assign new_n550_ = pi036 ^ pi037;
  assign new_n551_ = ~new_n552_ & ~pi039 & ~pi038;
  assign new_n552_ = ~new_n424_ | (~pi036 & pi037) | (pi036 & ~pi037);
  assign new_n553_ = new_n424_ & (~pi036 ^ pi037);
  assign new_n554_ = ~new_n556_ & ((~pi096 & (new_n445_ | ~new_n555_)) | ~new_n547_ | (~new_n445_ & ~new_n555_));
  assign new_n555_ = pi140 & pi097;
  assign new_n556_ = (~pi140 & pi096 & ~new_n551_) | (pi009 & ~new_n549_ & ~new_n550_);
  assign new_n557_ = ~new_n559_ & ((~pi097 & (new_n445_ | ~new_n558_)) | ~new_n547_ | (~new_n445_ & ~new_n558_));
  assign new_n558_ = pi140 & pi098;
  assign new_n559_ = (~pi140 & pi097 & ~new_n551_) | (pi010 & ~new_n549_ & ~new_n550_);
  assign new_n560_ = ~new_n562_ & ((~pi098 & (new_n445_ | ~new_n561_)) | ~new_n547_ | (~new_n445_ & ~new_n561_));
  assign new_n561_ = pi140 & pi099;
  assign new_n562_ = (~pi140 & pi098 & ~new_n551_) | (pi011 & ~new_n549_ & ~new_n550_);
  assign new_n563_ = ~new_n565_ & ((~pi099 & (new_n445_ | ~new_n564_)) | ~new_n547_ | (~new_n445_ & ~new_n564_));
  assign new_n564_ = pi140 & pi100;
  assign new_n565_ = (~pi140 & pi099 & ~new_n551_) | (pi012 & ~new_n549_ & ~new_n550_);
  assign new_n566_ = ~new_n568_ & ((~pi100 & (new_n445_ | ~new_n567_)) | ~new_n547_ | (~new_n445_ & ~new_n567_));
  assign new_n567_ = pi140 & pi101;
  assign new_n568_ = (~pi140 & pi100 & ~new_n551_) | (pi013 & ~new_n549_ & ~new_n550_);
  assign new_n569_ = ~new_n571_ & ((~pi101 & (new_n445_ | ~new_n570_)) | ~new_n547_ | (~new_n445_ & ~new_n570_));
  assign new_n570_ = pi140 & pi102;
  assign new_n571_ = (~pi140 & pi101 & ~new_n551_) | (pi014 & ~new_n549_ & ~new_n550_);
  assign new_n572_ = ~pi015 | pi039 | pi038;
  assign new_n573_ = ~pi040 | ~new_n424_ | pi042;
  assign new_n574_ = ~pi102 | pi042;
  assign new_n575_ = (~pi038 & ~new_n440_ & ~new_n550_) | (pi140 & ~new_n445_);
  assign new_n576_ = ~pi040 | ~new_n587_ | pi042;
  assign new_n577_ = new_n585_ | ~pi139 | ~pi104;
  assign new_n578_ = ~new_n593_ | (pi058 & ~new_n591_) | (pi059 & ~new_n592_);
  assign new_n579_ = ~pi103 | pi042;
  assign new_n580_ = ~new_n583_ & (~pi058 | ~new_n581_) & (~pi059 | ~new_n582_);
  assign new_n581_ = ~new_n590_ | pi060 | pi059;
  assign new_n582_ = pi060 | pi062 | pi061;
  assign new_n583_ = ~new_n584_ | ~pi139 | (pi062 & pi061);
  assign new_n584_ = ~new_n585_ & ~new_n586_ & (~pi062 | ~pi060);
  assign new_n585_ = ~pi136 & ~new_n804_;
  assign new_n586_ = ~new_n588_ | ~new_n587_ | (pi061 & pi060);
  assign new_n587_ = ~new_n788_ | (pi058 & ~pi048) | (pi059 & ~pi049);
  assign new_n588_ = ~new_n589_ | pi062 | pi061;
  assign new_n589_ = ~pi058 & ~pi060 & ~pi059;
  assign new_n590_ = ~pi062 & ~pi061;
  assign new_n591_ = ~new_n595_ & ~pi060 & ~pi059;
  assign new_n592_ = ~pi060 & ~pi062 & ~pi061;
  assign new_n593_ = ~new_n594_ & (pi059 | pi058 | ~new_n592_);
  assign new_n594_ = (pi061 & pi062) | (pi060 & (pi061 | pi062));
  assign new_n595_ = pi062 | pi061;
  assign new_n596_ = new_n585_ | ~pi139 | ~pi105;
  assign new_n597_ = ~pi104 | pi042;
  assign new_n598_ = new_n585_ | ~pi139 | ~pi106;
  assign new_n599_ = ~pi105 | pi042;
  assign new_n600_ = new_n585_ | ~pi139 | ~pi107;
  assign new_n601_ = ~pi106 | pi042;
  assign new_n602_ = new_n585_ | ~pi139 | ~pi108;
  assign new_n603_ = ~pi107 | pi042;
  assign new_n604_ = new_n585_ | ~pi139 | ~pi109;
  assign new_n605_ = ~pi108 | pi042;
  assign new_n606_ = new_n585_ | ~pi139 | ~pi110;
  assign new_n607_ = ~pi109 | pi042;
  assign new_n608_ = new_n585_ | ~pi139 | ~pi111;
  assign new_n609_ = ~pi110 | pi042;
  assign new_n610_ = new_n585_ | ~pi139 | ~pi112;
  assign new_n611_ = ~pi111 | pi042;
  assign new_n612_ = new_n585_ | ~pi139 | ~pi113;
  assign new_n613_ = ~pi112 | pi042;
  assign new_n614_ = new_n585_ | ~pi139 | ~pi114;
  assign new_n615_ = ~pi113 | pi042;
  assign new_n616_ = new_n585_ | ~pi139 | ~pi115;
  assign new_n617_ = ~pi114 | pi042;
  assign new_n618_ = new_n585_ | ~pi139 | ~pi116;
  assign new_n619_ = ~pi115 | pi042;
  assign new_n620_ = new_n585_ | ~pi139 | ~pi117;
  assign new_n621_ = ~pi116 | pi042;
  assign new_n622_ = new_n585_ | ~pi139 | ~pi118;
  assign new_n623_ = ~pi117 | pi042;
  assign new_n624_ = new_n585_ | ~pi139 | ~pi119;
  assign new_n625_ = ~pi118 | pi042;
  assign new_n626_ = new_n585_ | ~pi139 | ~pi120;
  assign new_n627_ = ~pi119 | pi042;
  assign new_n628_ = new_n585_ | ~pi139 | ~pi121;
  assign new_n629_ = ~pi120 | pi042;
  assign new_n630_ = new_n585_ | ~pi139 | ~pi122;
  assign new_n631_ = ~pi121 | pi042;
  assign new_n632_ = new_n585_ | ~pi139 | ~pi123;
  assign new_n633_ = ~pi122 | pi042;
  assign new_n634_ = new_n585_ | ~pi139 | ~pi124;
  assign new_n635_ = ~pi123 | pi042;
  assign new_n636_ = new_n585_ | ~pi139 | ~pi125;
  assign new_n637_ = ~pi124 | pi042;
  assign new_n638_ = pi042 | ~pi040;
  assign new_n639_ = ~new_n587_ | ~pi139 | new_n585_;
  assign new_n640_ = (pi058 | ~new_n648_) & (~pi043 | ~new_n647_ | ~new_n592_);
  assign new_n641_ = ~pi125 | pi042;
  assign new_n642_ = ~new_n643_ & (~pi058 | ~new_n581_) & (~pi059 | ~new_n582_);
  assign new_n643_ = ~new_n644_ | ~pi139 | new_n585_;
  assign new_n644_ = new_n587_ & ~new_n645_ & (~pi062 | ~pi061);
  assign new_n645_ = ~new_n646_ | (~pi059 & ~pi058 & ~new_n582_);
  assign new_n646_ = ~pi060 | (~pi061 & ~pi062);
  assign new_n647_ = ~pi059 & pi058;
  assign new_n648_ = pi059 ? (~new_n582_ & pi044) : ~new_n649_;
  assign new_n649_ = ~new_n651_ & (((~pi045 | ~new_n590_) & (~pi047 | pi060 | ~new_n650_)) | (~pi060 & (~pi047 | ~new_n650_)));
  assign new_n650_ = pi062 & ~pi061;
  assign new_n651_ = ~pi062 & ~new_n652_;
  assign new_n652_ = ~pi046 | ~pi061 | pi060;
  assign new_n653_ = ~new_n654_ | (pi140 & pi126 & ~new_n445_);
  assign new_n654_ = pi040 & ~pi042 & (pi039 | ~new_n424_);
  assign new_n655_ = ~new_n445_ & pi140 & ~pi126;
  assign new_n656_ = ~pi042 & ~new_n657_ & (~new_n424_ | pi039);
  assign new_n657_ = pi140 & ~new_n658_;
  assign new_n658_ = new_n445_ | pi127 | pi126;
  assign new_n659_ = ~new_n663_ & ~pi126 & ~new_n445_;
  assign new_n660_ = ~pi042 & ~new_n661_ & (~new_n424_ | pi039);
  assign new_n661_ = ~new_n662_ & pi140 & ~pi128;
  assign new_n662_ = new_n445_ | ~pi127 | pi126;
  assign new_n663_ = ~pi140 | ~pi127;
  assign new_n664_ = ~new_n668_ & (~new_n665_ | ~new_n666_ | ~new_n440_) & (~pi129 | ~pi039 | ~new_n667_);
  assign new_n665_ = ~new_n445_ & pi127 & ~pi126;
  assign new_n666_ = pi128 & pi140 & ~pi129;
  assign new_n667_ = ~new_n672_ | pi126 | new_n445_;
  assign new_n668_ = ~new_n669_ & ((pi129 & ~new_n424_) | ((pi129 | new_n424_) & (pi038 | ~new_n550_)));
  assign new_n669_ = new_n424_ ? pi039 : (~new_n670_ & ~new_n671_);
  assign new_n670_ = pi126 | new_n445_;
  assign new_n671_ = ~pi127 | ~pi140 | ~pi128;
  assign new_n672_ = pi127 & pi140 & pi128;
  assign new_n673_ = ~new_n683_ | ~pi040 | ~new_n682_;
  assign new_n674_ = pi042 | pi126 | new_n445_;
  assign new_n675_ = new_n424_ & ~pi039;
  assign new_n676_ = ~pi130 | pi042;
  assign new_n677_ = (~new_n445_ & ~new_n680_ & ~new_n681_) | (new_n424_ & ~pi039);
  assign new_n678_ = ~new_n679_ | ~new_n424_ | pi042;
  assign new_n679_ = pi038 & pi040 & ~pi039;
  assign new_n680_ = ~pi127 | pi126;
  assign new_n681_ = ~pi128 | ~pi140 | pi129;
  assign new_n682_ = pi128 & pi127;
  assign new_n683_ = ~pi129 & pi140 & ~pi130;
  assign new_n684_ = ~new_n692_ | ~pi040 | ~new_n691_;
  assign new_n685_ = ~pi131 | pi042;
  assign new_n686_ = (~new_n445_ & ~new_n689_ & ~new_n690_) | (new_n424_ & ~pi039);
  assign new_n687_ = ~new_n688_ | ~new_n424_ | pi042;
  assign new_n688_ = ~pi038 & pi040 & ~pi039;
  assign new_n689_ = pi126 | ~pi128 | ~pi127;
  assign new_n690_ = pi129 | ~pi140 | pi130;
  assign new_n691_ = pi127 & ~pi129 & pi128;
  assign new_n692_ = ~pi130 & pi140 & ~pi131;
  assign new_n693_ = pi057 | pi042;
  assign new_n694_ = (~pi132 & ~new_n697_) | (~new_n585_ & new_n587_ & ~new_n696_);
  assign new_n695_ = ~new_n424_ | pi042;
  assign new_n696_ = ~pi139 | ~pi132;
  assign new_n697_ = new_n587_ & pi139 & ~new_n585_;
  assign new_n698_ = ~new_n702_ & ~new_n585_ & new_n587_;
  assign new_n699_ = ~new_n700_ & ~pi042 & ~pi057;
  assign new_n700_ = (new_n424_ & ~pi039) | (~new_n585_ & new_n587_ & ~new_n701_);
  assign new_n701_ = pi132 | ~pi139 | pi133;
  assign new_n702_ = ~pi139 | pi132;
  assign new_n703_ = ~new_n708_ & ~new_n585_ & new_n587_;
  assign new_n704_ = ~new_n705_ & ~pi042 & ~pi057;
  assign new_n705_ = (new_n587_ & ~new_n706_ & ~new_n707_) | (new_n424_ & ~pi039);
  assign new_n706_ = pi132 | new_n585_;
  assign new_n707_ = ~pi133 | ~pi139 | pi134;
  assign new_n708_ = pi132 | ~pi139 | ~pi133;
  assign new_n709_ = ~new_n718_ | ~pi040 | ~new_n717_;
  assign new_n710_ = pi042 | new_n585_ | ~new_n587_;
  assign new_n711_ = pi042 | ~pi135 | pi057;
  assign new_n712_ = (new_n587_ & ~new_n706_ & ~new_n716_) | (new_n424_ & ~pi039);
  assign new_n713_ = ~new_n714_ | ~new_n424_ | pi042;
  assign new_n714_ = pi040 & ~new_n715_;
  assign new_n715_ = pi039 | (pi038 & (pi036 ^ pi037));
  assign new_n716_ = ~pi133 | ~pi139 | ~pi134;
  assign new_n717_ = ~pi057 & pi133 & ~pi132;
  assign new_n718_ = pi134 & pi139 & ~pi135;
  assign new_n719_ = ~new_n726_ | ~new_n724_ | ~new_n725_;
  assign new_n720_ = pi042 | ~pi136 | pi057;
  assign new_n721_ = (new_n587_ & ~new_n722_ & ~new_n723_) | (new_n424_ & ~pi039);
  assign new_n722_ = new_n585_ | ~pi133 | pi132;
  assign new_n723_ = ~pi134 | ~pi139 | pi135;
  assign new_n724_ = ~pi057 & ~new_n585_;
  assign new_n725_ = ~pi132 & pi134 & pi133;
  assign new_n726_ = ~pi135 & pi139 & ~pi136;
  assign new_n727_ = ~new_n728_ | (pi137 & pi064);
  assign new_n728_ = pi040 & ~new_n445_ & ~pi042;
  assign new_n729_ = ~new_n742_ | pi042 | ~pi040;
  assign new_n730_ = ~new_n587_ | pi057 | new_n585_;
  assign new_n731_ = pi042 | ~pi138 | pi057;
  assign new_n732_ = ~new_n736_ & ((pi058 & ~new_n735_) | ((~pi058 | ~new_n735_) & (~new_n733_ | ~new_n734_)));
  assign new_n733_ = ~pi060 & ~pi059;
  assign new_n734_ = (~pi046 & ~pi062) | (~pi061 & (~pi047 | ~pi062));
  assign new_n735_ = ~new_n592_ | pi059 | ~pi043;
  assign new_n736_ = ~new_n739_ | (~pi058 & ~pi045 & ~new_n737_) | (pi059 & ~new_n738_);
  assign new_n737_ = pi059 | pi062 | pi061;
  assign new_n738_ = ~new_n595_ & ~pi060 & pi044;
  assign new_n739_ = ~new_n740_ & pi142 & pi139;
  assign new_n740_ = ~new_n741_ | ~new_n587_ | (pi062 & pi061);
  assign new_n741_ = ~new_n585_ & (~pi060 | (~pi061 & ~pi062));
  assign new_n742_ = ~pi138 & pi142 & pi139;
  assign new_n743_ = ~new_n691_ | ~pi040 | ~new_n744_;
  assign new_n744_ = pi063 & ~pi042;
  assign new_n745_ = ~pi040 | new_n445_ | pi042;
  assign new_n746_ = ~new_n789_ | ~pi142 | (pi058 & ~pi048);
  assign new_n747_ = ~pi040 | pi042 | (~new_n587_ & new_n746_);
  assign new_n748_ = (~pi106 & (~pi037 | ~pi114)) | (pi037 & ~pi114);
  assign new_n749_ = (~pi106 & (pi037 | ~pi114)) | (~pi037 & ~pi114);
  assign new_n750_ = ~pi122 & ~pi038;
  assign new_n751_ = (~pi105 & (~pi037 | ~pi113)) | (pi037 & ~pi113);
  assign new_n752_ = (~pi105 & (pi037 | ~pi113)) | (~pi037 & ~pi113);
  assign new_n753_ = ~pi121 & ~pi038;
  assign new_n754_ = (~pi104 & (~pi037 | ~pi112)) | (pi037 & ~pi112);
  assign new_n755_ = (~pi104 & (pi037 | ~pi112)) | (~pi037 & ~pi112);
  assign new_n756_ = ~pi120 & ~pi038;
  assign new_n757_ = (~pi103 & (~pi037 | ~pi111)) | (pi037 & ~pi111);
  assign new_n758_ = (~pi103 & (pi037 | ~pi111)) | (~pi037 & ~pi111);
  assign new_n759_ = ~pi119 & ~pi038;
  assign new_n760_ = ~pi038 | (~pi107 & (~pi036 ^ pi037));
  assign new_n761_ = ~pi038 | (~pi108 & (~pi036 ^ pi037));
  assign new_n762_ = ~pi038 | (~pi109 & (~pi036 ^ pi037));
  assign new_n763_ = ~pi038 | (~pi110 & (~pi036 ^ pi037));
  assign new_n764_ = ~pi038 | (~pi111 & (~pi036 ^ pi037));
  assign new_n765_ = ~pi038 | (~pi112 & (~pi036 ^ pi037));
  assign new_n766_ = ~pi038 | (~pi113 & (~pi036 ^ pi037));
  assign new_n767_ = ~pi038 | (~pi114 & (~pi036 ^ pi037));
  assign new_n768_ = ~pi039 & ~pi139 & pi058;
  assign new_n769_ = ~pi039 & ~pi139 & pi059;
  assign new_n770_ = ~pi039 & ~pi139 & pi060;
  assign new_n771_ = ~pi039 & ~pi139 & pi061;
  assign new_n772_ = ~pi039 & ~pi139 & pi062;
  assign new_n773_ = ~pi129 & ~pi131 & ~pi130;
  assign new_n774_ = pi056 ^ pi137;
  assign new_n775_ = ~new_n773_ | ~pi128 | ~pi127;
  assign new_n776_ = pi058 & ~pi139 & pi063;
  assign new_n777_ = pi059 & ~pi139 & pi063;
  assign new_n778_ = pi060 & ~pi139 & pi063;
  assign new_n779_ = pi061 & ~pi139 & pi063;
  assign new_n780_ = pi062 & ~pi139 & pi063;
  assign new_n781_ = pi140 & pi058;
  assign new_n782_ = pi140 & pi059;
  assign new_n783_ = pi140 & pi060;
  assign new_n784_ = pi140 & pi061;
  assign new_n785_ = pi140 & pi062;
  assign new_n786_ = ~new_n787_ | ~pi127 | ~pi126;
  assign new_n787_ = ~pi129 & pi128;
  assign new_n788_ = (pi052 | ~pi062) & (pi050 | ~pi060) & (pi051 | ~pi061);
  assign new_n789_ = ~new_n790_ & (~pi059 | pi049) & (~pi060 | pi050);
  assign new_n790_ = ~new_n791_ | (pi061 & ~pi051) | (pi062 & ~pi052);
  assign new_n791_ = pi136 | ~new_n792_;
  assign new_n792_ = pi133 & ~pi135 & pi134;
  assign new_n793_ = ~new_n801_ & pi134 & pi133;
  assign new_n794_ = ~new_n796_ & (~new_n795_ | ((~pi060 | pi050) & (~pi061 | pi051)));
  assign new_n795_ = ~new_n800_ | ~pi134 | ~pi133;
  assign new_n796_ = ~new_n797_ & (~pi142 | ~new_n795_ | (~pi052 & pi062));
  assign new_n797_ = ~new_n798_ & ~pi136 & ~pi135;
  assign new_n798_ = ~new_n799_ | ~pi132 | pi057;
  assign new_n799_ = pi134 & pi133;
  assign new_n800_ = ~pi136 & ~pi135;
  assign new_n801_ = pi136 | pi135;
  assign new_n802_ = pi058 | pi060 | pi059;
  assign new_n803_ = ~new_n787_ | ~pi127 | pi126;
  assign new_n804_ = ~pi133 | pi135 | ~pi134;
  assign po005 = pi123;
  assign po006 = pi124;
  assign po024 = pi141;
  assign po050 = pi139;
endmodule


