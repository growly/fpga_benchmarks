// Benchmark "C2670.iscas" written by ABC on Thu Mar 19 13:02:35 2020

module C2670_iscas  ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139;
  wire new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n441_, new_n449_, new_n451_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n491_, new_n492_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n518_, new_n519_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n765_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n834_, new_n836_, new_n838_, new_n840_, new_n842_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_,
    new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_,
    new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_,
    new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_,
    new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_,
    new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_,
    new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_,
    new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_,
    new_n1185_, new_n1186_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_,
    new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_,
    new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_,
    new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_,
    new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_,
    new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_,
    new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_,
    new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_,
    new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_,
    new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_,
    new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_,
    new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1322_, new_n1323_, new_n1324_, new_n1325_,
    new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_,
    new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_,
    new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_,
    new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_,
    new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_,
    new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_,
    new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_,
    new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_,
    new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_,
    new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_,
    new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_,
    new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_,
    new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_,
    new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_,
    new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_,
    new_n1416_, new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_,
    new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_,
    new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_,
    new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_,
    new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_,
    new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_,
    new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_,
    new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_,
    new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_,
    new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_,
    new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_,
    new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_,
    new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_,
    new_n1497_, new_n1498_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_,
    new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_,
    new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_,
    new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1534_,
    new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1548_, new_n1549_,
    new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_,
    new_n1564_;
  assign new_n374_ = ~pi232;
  assign new_n375_ = ~pi231;
  assign new_n376_ = ~pi230;
  assign new_n377_ = ~pi229;
  assign new_n378_ = ~pi228;
  assign new_n379_ = ~pi227;
  assign new_n380_ = ~pi226;
  assign new_n381_ = ~pi225;
  assign new_n382_ = ~pi224;
  assign new_n383_ = ~pi223;
  assign new_n384_ = pi221;
  assign new_n385_ = pi221;
  assign new_n386_ = pi220;
  assign new_n387_ = pi220;
  assign new_n388_ = ~pi219;
  assign new_n389_ = pi219;
  assign new_n390_ = ~pi218;
  assign new_n391_ = pi218;
  assign new_n392_ = ~pi217;
  assign new_n393_ = pi217;
  assign new_n394_ = ~pi216;
  assign new_n395_ = pi216;
  assign new_n396_ = ~pi215;
  assign new_n397_ = pi215;
  assign new_n398_ = ~pi214;
  assign new_n399_ = pi214;
  assign new_n400_ = pi214 & pi215 & pi217 & pi216;
  assign new_n401_ = ~pi213;
  assign new_n402_ = pi213;
  assign po083 = pi212;
  assign po082 = pi212;
  assign po081 = pi212;
  assign new_n406_ = ~pi211;
  assign new_n407_ = pi211;
  assign new_n408_ = ~pi210;
  assign new_n409_ = pi210;
  assign new_n410_ = ~pi209;
  assign new_n411_ = pi209;
  assign new_n412_ = ~pi208;
  assign new_n413_ = pi208;
  assign new_n414_ = ~pi207;
  assign new_n415_ = pi207;
  assign new_n416_ = ~pi206;
  assign new_n417_ = pi206;
  assign new_n418_ = ~pi205;
  assign new_n419_ = pi205;
  assign new_n420_ = ~pi204;
  assign new_n421_ = pi204;
  assign new_n422_ = ~pi203;
  assign new_n423_ = pi203;
  assign new_n424_ = ~pi202;
  assign new_n425_ = ~pi201;
  assign new_n426_ = pi201;
  assign new_n427_ = ~pi200;
  assign new_n428_ = pi200;
  assign po080 = pi199;
  assign po079 = pi199;
  assign new_n431_ = ~pi198;
  assign new_n432_ = ~pi197;
  assign new_n433_ = pi196;
  assign new_n434_ = pi195;
  assign new_n435_ = pi195;
  assign new_n436_ = ~pi193;
  assign new_n437_ = pi192;
  assign new_n438_ = pi192;
  assign po078 = pi190;
  assign po077 = pi190;
  assign new_n441_ = pi190;
  assign po076 = pi190;
  assign po085 = ~pi105;
  assign po089 = ~pi095;
  assign po091 = ~pi085;
  assign po087 = ~pi075;
  assign po086 = ~pi063;
  assign po088 = ~pi052;
  assign new_n449_ = pi052 & pi085 & pi095 & pi042;
  assign po090 = ~pi042;
  assign new_n451_ = pi031 & pi075 & pi105 & pi063;
  assign po084 = ~pi031;
  assign new_n453_ = pi028 & pi028;
  assign new_n454_ = pi022;
  assign new_n455_ = pi022;
  assign new_n456_ = pi011;
  assign new_n457_ = pi011;
  assign new_n458_ = pi008 & pi198;
  assign new_n459_ = pi007;
  assign new_n460_ = pi007;
  assign new_n461_ = pi006 & pi196;
  assign new_n462_ = pi196 & pi001 & pi010;
  assign new_n463_ = pi000 & pi002;
  assign new_n464_ = ~new_n402_ | ~new_n374_;
  assign new_n465_ = ~new_n423_ | ~new_n375_;
  assign new_n466_ = ~pi230 | ~new_n377_;
  assign new_n467_ = ~pi229 | ~new_n376_;
  assign new_n468_ = ~pi228 | ~new_n379_;
  assign new_n469_ = ~pi227 | ~new_n378_;
  assign new_n470_ = ~pi226 | ~new_n381_;
  assign new_n471_ = ~pi225 | ~new_n380_;
  assign new_n472_ = ~pi224 | ~new_n383_;
  assign new_n473_ = ~pi223 | ~new_n382_;
  assign new_n474_ = pi222 & new_n461_;
  assign new_n475_ = ~new_n384_;
  assign new_n476_ = new_n387_ & new_n385_;
  assign new_n477_ = ~new_n385_;
  assign new_n478_ = ~new_n386_;
  assign new_n479_ = ~new_n387_;
  assign new_n480_ = ~new_n389_;
  assign new_n481_ = ~new_n391_;
  assign new_n482_ = new_n392_;
  assign new_n483_ = ~new_n393_;
  assign new_n484_ = new_n394_;
  assign new_n485_ = ~new_n395_;
  assign new_n486_ = new_n396_;
  assign new_n487_ = ~new_n397_;
  assign new_n488_ = new_n398_;
  assign new_n489_ = ~new_n399_;
  assign po092 = ~new_n400_;
  assign new_n491_ = new_n401_;
  assign new_n492_ = ~new_n402_;
  assign new_n493_ = new_n406_;
  assign new_n494_ = ~new_n407_;
  assign new_n495_ = new_n408_;
  assign new_n496_ = ~new_n409_;
  assign new_n497_ = new_n410_;
  assign new_n498_ = ~new_n411_;
  assign new_n499_ = new_n412_;
  assign new_n500_ = ~new_n413_;
  assign new_n501_ = new_n414_;
  assign new_n502_ = ~new_n415_;
  assign new_n503_ = new_n416_;
  assign new_n504_ = ~new_n417_;
  assign new_n505_ = new_n418_;
  assign new_n506_ = ~new_n419_;
  assign new_n507_ = new_n420_;
  assign new_n508_ = ~new_n421_;
  assign new_n509_ = new_n422_;
  assign new_n510_ = ~new_n423_;
  assign new_n511_ = new_n425_;
  assign new_n512_ = ~new_n426_;
  assign new_n513_ = new_n427_;
  assign new_n514_ = ~new_n428_;
  assign new_n515_ = ~new_n434_;
  assign new_n516_ = ~new_n435_;
  assign po097 = ~pi194 | ~new_n461_;
  assign new_n518_ = ~new_n437_;
  assign new_n519_ = ~new_n438_;
  assign po094 = new_n441_;
  assign new_n521_ = new_n384_ & pi093 & new_n386_;
  assign new_n522_ = new_n384_ & pi092 & new_n386_;
  assign new_n523_ = new_n384_ & pi091 & new_n386_;
  assign new_n524_ = new_n384_ & pi090 & new_n386_;
  assign new_n525_ = new_n385_ & pi089 & new_n387_;
  assign new_n526_ = new_n385_ & pi088 & new_n387_;
  assign new_n527_ = new_n385_ & pi087 & new_n387_;
  assign new_n528_ = new_n385_ & pi086 & new_n387_;
  assign new_n529_ = new_n384_ & pi084 & new_n386_;
  assign po095 = pi073 & new_n441_;
  assign new_n531_ = new_n435_ & pi061 & new_n438_;
  assign new_n532_ = new_n435_ & pi060 & new_n438_;
  assign new_n533_ = new_n435_ & pi059 & new_n438_;
  assign new_n534_ = new_n435_ & pi058 & new_n438_;
  assign new_n535_ = new_n434_ & pi057 & new_n437_;
  assign new_n536_ = new_n434_ & pi056 & new_n437_;
  assign new_n537_ = new_n434_ & pi055 & new_n437_;
  assign new_n538_ = new_n434_ & pi054 & new_n437_;
  assign new_n539_ = new_n434_ & pi053 & new_n437_;
  assign new_n540_ = new_n435_ & pi051 & new_n438_;
  assign new_n541_ = new_n449_ & new_n451_;
  assign new_n542_ = ~new_n449_;
  assign new_n543_ = ~new_n451_;
  assign new_n544_ = ~new_n453_;
  assign new_n545_ = ~new_n454_;
  assign new_n546_ = ~new_n455_;
  assign new_n547_ = ~new_n456_;
  assign new_n548_ = ~new_n457_;
  assign new_n549_ = pi008 & new_n431_;
  assign new_n550_ = new_n459_;
  assign new_n551_ = new_n459_;
  assign new_n552_ = new_n460_;
  assign new_n553_ = new_n460_;
  assign po096 = ~new_n461_;
  assign po093 = ~new_n462_;
  assign new_n556_ = ~new_n463_;
  assign new_n557_ = ~pi232 | ~new_n492_;
  assign new_n558_ = ~pi231 | ~new_n510_;
  assign new_n559_ = ~new_n466_ | ~new_n467_;
  assign new_n560_ = ~new_n468_ | ~new_n469_;
  assign new_n561_ = ~new_n470_ | ~new_n471_;
  assign new_n562_ = ~new_n472_ | ~new_n473_;
  assign new_n563_ = pi222 & new_n543_;
  assign po098 = ~new_n474_;
  assign new_n565_ = new_n479_ & new_n385_;
  assign new_n566_ = new_n479_ & new_n477_;
  assign new_n567_ = new_n387_ & new_n477_;
  assign new_n568_ = ~new_n389_ | ~new_n481_;
  assign new_n569_ = ~new_n391_ | ~new_n480_;
  assign new_n570_ = ~new_n482_;
  assign new_n571_ = ~new_n393_ | ~new_n485_;
  assign new_n572_ = ~new_n484_;
  assign new_n573_ = ~new_n395_ | ~new_n483_;
  assign new_n574_ = ~new_n486_;
  assign new_n575_ = ~new_n397_ | ~new_n489_;
  assign new_n576_ = ~new_n488_;
  assign new_n577_ = ~new_n399_ | ~new_n487_;
  assign new_n578_ = ~new_n491_;
  assign new_n579_ = ~new_n493_;
  assign new_n580_ = ~new_n407_ | ~new_n496_;
  assign new_n581_ = ~new_n495_;
  assign new_n582_ = ~new_n409_ | ~new_n494_;
  assign new_n583_ = ~new_n497_;
  assign new_n584_ = ~new_n411_ | ~new_n500_;
  assign new_n585_ = ~new_n499_;
  assign new_n586_ = ~new_n413_ | ~new_n498_;
  assign new_n587_ = ~new_n501_;
  assign new_n588_ = ~new_n415_ | ~new_n504_;
  assign new_n589_ = ~new_n503_;
  assign new_n590_ = ~new_n417_ | ~new_n502_;
  assign new_n591_ = ~new_n505_;
  assign new_n592_ = ~new_n419_ | ~new_n508_;
  assign new_n593_ = ~new_n507_;
  assign new_n594_ = ~new_n421_ | ~new_n506_;
  assign new_n595_ = ~new_n509_;
  assign new_n596_ = ~new_n511_;
  assign new_n597_ = ~new_n426_ | ~new_n514_;
  assign new_n598_ = ~new_n513_;
  assign new_n599_ = ~new_n428_ | ~new_n512_;
  assign new_n600_ = new_n518_ & new_n434_;
  assign new_n601_ = pi194 & new_n542_;
  assign new_n602_ = new_n475_ & pi113 & new_n478_;
  assign new_n603_ = new_n475_ & pi112 & new_n478_;
  assign new_n604_ = new_n475_ & pi111 & new_n478_;
  assign new_n605_ = new_n475_ & pi110 & new_n478_;
  assign new_n606_ = new_n477_ & pi109 & new_n479_;
  assign new_n607_ = new_n477_ & pi108 & new_n479_;
  assign new_n608_ = new_n477_ & pi107 & new_n479_;
  assign new_n609_ = new_n477_ & pi106 & new_n479_;
  assign new_n610_ = new_n475_ & pi104 & new_n478_;
  assign new_n611_ = new_n384_ & pi103 & new_n478_;
  assign new_n612_ = new_n384_ & pi102 & new_n478_;
  assign new_n613_ = new_n384_ & pi101 & new_n478_;
  assign new_n614_ = new_n384_ & pi100 & new_n478_;
  assign new_n615_ = new_n385_ & pi099 & new_n479_;
  assign new_n616_ = new_n385_ & pi098 & new_n479_;
  assign new_n617_ = new_n385_ & pi097 & new_n479_;
  assign new_n618_ = new_n385_ & pi096 & new_n479_;
  assign new_n619_ = new_n384_ & pi094 & new_n478_;
  assign new_n620_ = new_n475_ & pi083 & new_n386_;
  assign new_n621_ = new_n475_ & pi082 & new_n386_;
  assign new_n622_ = new_n475_ & pi081 & new_n386_;
  assign new_n623_ = new_n475_ & pi080 & new_n386_;
  assign new_n624_ = new_n477_ & pi079 & new_n387_;
  assign new_n625_ = new_n477_ & pi078 & new_n387_;
  assign new_n626_ = new_n477_ & pi077 & new_n387_;
  assign new_n627_ = new_n477_ & pi076 & new_n387_;
  assign new_n628_ = new_n475_ & pi074 & new_n386_;
  assign new_n629_ = new_n516_ & pi072 & new_n519_;
  assign new_n630_ = new_n516_ & pi071 & new_n519_;
  assign new_n631_ = new_n516_ & pi070 & new_n519_;
  assign new_n632_ = new_n516_ & pi069 & new_n519_;
  assign new_n633_ = new_n515_ & pi068 & new_n518_;
  assign new_n634_ = new_n515_ & pi067 & new_n518_;
  assign new_n635_ = new_n515_ & pi066 & new_n518_;
  assign new_n636_ = new_n515_ & pi065 & new_n518_;
  assign new_n637_ = new_n515_ & pi064 & new_n518_;
  assign new_n638_ = new_n516_ & pi062 & new_n519_;
  assign new_n639_ = new_n435_ & pi050 & new_n519_;
  assign new_n640_ = new_n435_ & pi049 & new_n519_;
  assign new_n641_ = new_n435_ & pi048 & new_n519_;
  assign new_n642_ = new_n435_ & pi047 & new_n519_;
  assign new_n643_ = new_n434_ & pi046 & new_n518_;
  assign new_n644_ = new_n434_ & pi045 & new_n518_;
  assign new_n645_ = new_n434_ & pi044 & new_n518_;
  assign new_n646_ = new_n434_ & pi043 & new_n518_;
  assign po100 = ~new_n541_;
  assign po099 = new_n541_;
  assign new_n649_ = new_n435_ & pi041 & new_n519_;
  assign new_n650_ = new_n516_ & pi040 & new_n438_;
  assign new_n651_ = new_n516_ & pi039 & new_n438_;
  assign new_n652_ = new_n516_ & pi038 & new_n438_;
  assign new_n653_ = new_n516_ & pi037 & new_n438_;
  assign new_n654_ = new_n515_ & pi036 & new_n437_;
  assign new_n655_ = new_n515_ & pi035 & new_n437_;
  assign new_n656_ = new_n515_ & pi034 & new_n437_;
  assign new_n657_ = new_n515_ & pi033 & new_n437_;
  assign new_n658_ = new_n515_ & pi032 & new_n437_;
  assign new_n659_ = new_n516_ & pi030 & new_n438_;
  assign new_n660_ = pi026 & new_n545_;
  assign new_n661_ = pi025 & new_n545_;
  assign new_n662_ = pi024 & new_n546_;
  assign new_n663_ = pi023 & new_n546_;
  assign new_n664_ = pi021 & new_n545_;
  assign new_n665_ = pi020 & new_n545_;
  assign new_n666_ = pi019 & new_n546_;
  assign new_n667_ = pi018 & new_n546_;
  assign new_n668_ = pi017 & new_n547_;
  assign new_n669_ = pi016 & new_n547_;
  assign new_n670_ = pi015 & new_n547_;
  assign new_n671_ = pi014 & new_n547_;
  assign new_n672_ = pi013 & new_n548_;
  assign new_n673_ = pi012 & new_n548_;
  assign new_n674_ = new_n549_ | new_n458_;
  assign new_n675_ = pi005 & new_n547_;
  assign new_n676_ = pi004 & new_n548_;
  assign new_n677_ = pi003 & new_n548_;
  assign new_n678_ = ~new_n557_ | ~new_n464_;
  assign new_n679_ = ~new_n558_ | ~new_n465_;
  assign new_n680_ = ~new_n559_;
  assign new_n681_ = new_n560_;
  assign new_n682_ = new_n560_;
  assign new_n683_ = ~new_n561_;
  assign new_n684_ = ~new_n562_;
  assign new_n685_ = ~new_n563_;
  assign new_n686_ = new_n476_ | new_n565_ | new_n566_ | new_n567_;
  assign new_n687_ = ~new_n569_ | ~new_n568_;
  assign new_n688_ = ~new_n573_ | ~new_n571_;
  assign new_n689_ = ~new_n577_ | ~new_n575_;
  assign new_n690_ = ~new_n582_ | ~new_n580_;
  assign new_n691_ = ~new_n586_ | ~new_n584_;
  assign new_n692_ = ~new_n590_ | ~new_n588_;
  assign new_n693_ = ~new_n594_ | ~new_n592_;
  assign new_n694_ = ~new_n599_ | ~new_n597_;
  assign new_n695_ = ~new_n601_;
  assign new_n696_ = new_n521_ | new_n611_ | new_n602_ | new_n620_;
  assign new_n697_ = new_n522_ | new_n612_ | new_n603_ | new_n621_;
  assign new_n698_ = new_n523_ | new_n613_ | new_n604_ | new_n622_;
  assign new_n699_ = new_n524_ | new_n614_ | new_n605_ | new_n623_;
  assign new_n700_ = new_n525_ | new_n615_ | new_n606_ | new_n624_;
  assign new_n701_ = new_n526_ | new_n616_ | new_n607_ | new_n625_;
  assign new_n702_ = new_n527_ | new_n617_ | new_n608_ | new_n626_;
  assign new_n703_ = new_n528_ | new_n618_ | new_n609_ | new_n627_;
  assign new_n704_ = new_n529_ | new_n619_ | new_n610_ | new_n628_;
  assign new_n705_ = new_n531_ | new_n639_ | new_n629_ | new_n650_;
  assign new_n706_ = new_n532_ | new_n640_ | new_n630_ | new_n651_;
  assign new_n707_ = new_n533_ | new_n641_ | new_n631_ | new_n652_;
  assign new_n708_ = new_n534_ | new_n642_ | new_n632_ | new_n653_;
  assign new_n709_ = new_n535_ | new_n643_ | new_n633_ | new_n654_;
  assign new_n710_ = new_n536_ | new_n644_ | new_n634_ | new_n655_;
  assign new_n711_ = new_n537_ | new_n600_ | new_n635_ | new_n656_;
  assign new_n712_ = new_n538_ | new_n645_ | new_n636_ | new_n657_;
  assign new_n713_ = new_n539_ | new_n646_ | new_n637_ | new_n658_;
  assign new_n714_ = new_n540_ | new_n649_ | new_n638_ | new_n659_;
  assign new_n715_ = ~new_n678_;
  assign new_n716_ = ~new_n679_;
  assign new_n717_ = ~new_n694_ | ~new_n680_;
  assign new_n718_ = new_n681_ & new_n683_ & new_n684_;
  assign new_n719_ = ~new_n681_;
  assign new_n720_ = ~new_n682_;
  assign new_n721_ = new_n682_ & new_n561_ & new_n562_;
  assign new_n722_ = new_n685_ & new_n695_;
  assign new_n723_ = new_n686_;
  assign new_n724_ = ~new_n388_ | ~new_n686_;
  assign new_n725_ = ~new_n687_;
  assign new_n726_ = ~new_n390_ | ~new_n703_;
  assign new_n727_ = new_n688_;
  assign new_n728_ = new_n688_;
  assign new_n729_ = ~new_n689_;
  assign new_n730_ = ~new_n690_;
  assign new_n731_ = ~new_n691_;
  assign new_n732_ = new_n692_;
  assign new_n733_ = new_n692_;
  assign new_n734_ = ~new_n693_;
  assign new_n735_ = new_n700_ & new_n424_;
  assign new_n736_ = ~new_n694_;
  assign new_n737_ = new_n714_ & new_n431_;
  assign new_n738_ = new_n706_ & new_n431_;
  assign new_n739_ = new_n709_ & pi198;
  assign new_n740_ = new_n714_ & pi197;
  assign new_n741_ = new_n706_ & pi197;
  assign new_n742_ = new_n705_ & pi197;
  assign new_n743_ = ~new_n696_;
  assign new_n744_ = new_n697_;
  assign new_n745_ = new_n698_;
  assign new_n746_ = new_n698_;
  assign new_n747_ = new_n699_;
  assign po104 = ~new_n700_;
  assign new_n749_ = new_n700_;
  assign po102 = ~new_n701_;
  assign new_n751_ = ~new_n701_;
  assign new_n752_ = new_n701_;
  assign po103 = ~new_n702_;
  assign new_n754_ = new_n702_;
  assign new_n755_ = new_n703_;
  assign new_n756_ = new_n704_;
  assign new_n757_ = new_n705_;
  assign new_n758_ = ~new_n705_;
  assign new_n759_ = ~new_n706_;
  assign new_n760_ = ~new_n706_;
  assign new_n761_ = new_n707_;
  assign po107 = ~new_n708_;
  assign new_n763_ = new_n708_;
  assign po106 = ~new_n709_;
  assign new_n765_ = new_n709_;
  assign po105 = ~new_n710_;
  assign new_n767_ = new_n710_;
  assign new_n768_ = new_n711_;
  assign new_n769_ = new_n712_;
  assign new_n770_ = new_n713_;
  assign new_n771_ = ~new_n714_;
  assign new_n772_ = new_n714_;
  assign new_n773_ = new_n702_ & new_n454_;
  assign new_n774_ = new_n701_ & new_n454_;
  assign new_n775_ = new_n700_ & new_n454_;
  assign new_n776_ = new_n703_ & new_n454_;
  assign new_n777_ = new_n704_ & new_n455_;
  assign new_n778_ = new_n699_ & new_n455_;
  assign new_n779_ = new_n698_ & new_n455_;
  assign new_n780_ = new_n697_ & new_n455_;
  assign new_n781_ = new_n711_ & new_n456_;
  assign new_n782_ = new_n710_ & new_n456_;
  assign new_n783_ = new_n709_ & new_n456_;
  assign new_n784_ = new_n713_ & new_n456_;
  assign new_n785_ = new_n712_ & new_n456_;
  assign new_n786_ = new_n714_ & new_n457_;
  assign new_n787_ = new_n708_ & new_n457_;
  assign new_n788_ = new_n707_ & new_n457_;
  assign new_n789_ = new_n706_ & new_n457_;
  assign new_n790_ = new_n728_ & new_n689_ & new_n678_;
  assign new_n791_ = new_n727_ & new_n729_ & new_n715_;
  assign new_n792_ = new_n733_ & new_n693_ & new_n679_;
  assign new_n793_ = new_n732_ & new_n734_ & new_n716_;
  assign new_n794_ = ~new_n559_ | ~new_n736_;
  assign new_n795_ = new_n720_ & new_n684_ & new_n561_;
  assign new_n796_ = new_n719_ & new_n562_ & new_n683_;
  assign po101 = new_n722_;
  assign new_n798_ = new_n724_ & new_n686_;
  assign new_n799_ = ~new_n723_;
  assign new_n800_ = new_n388_ & new_n724_;
  assign new_n801_ = new_n390_ & new_n726_;
  assign new_n802_ = ~new_n727_;
  assign new_n803_ = ~new_n728_;
  assign new_n804_ = ~new_n690_ | ~new_n731_;
  assign new_n805_ = ~new_n691_ | ~new_n730_;
  assign new_n806_ = ~new_n732_;
  assign new_n807_ = ~new_n733_;
  assign new_n808_ = ~new_n735_;
  assign new_n809_ = new_n757_ & new_n431_;
  assign new_n810_ = new_n761_ & new_n431_;
  assign new_n811_ = new_n763_ & pi198;
  assign po108 = new_n432_ | new_n740_;
  assign new_n813_ = ~new_n436_ | ~new_n760_;
  assign new_n814_ = new_n556_ & new_n722_ & new_n433_ & pi191;
  assign new_n815_ = ~new_n756_ | ~new_n743_;
  assign new_n816_ = ~new_n744_;
  assign new_n817_ = ~new_n746_;
  assign new_n818_ = ~new_n747_;
  assign new_n819_ = ~new_n749_;
  assign new_n820_ = ~new_n752_;
  assign new_n821_ = ~new_n754_;
  assign new_n822_ = new_n726_ & new_n703_;
  assign new_n823_ = ~new_n755_;
  assign new_n824_ = ~new_n756_;
  assign new_n825_ = new_n757_;
  assign new_n826_ = new_n758_;
  assign new_n827_ = new_n758_;
  assign new_n828_ = new_n759_;
  assign new_n829_ = new_n759_;
  assign new_n830_ = new_n759_;
  assign new_n831_ = new_n759_;
  assign new_n832_ = ~new_n760_;
  assign po111 = new_n761_;
  assign new_n834_ = ~new_n761_;
  assign po112 = new_n763_;
  assign new_n836_ = ~new_n763_;
  assign po113 = new_n765_;
  assign new_n838_ = ~new_n765_;
  assign po114 = new_n767_;
  assign new_n840_ = ~new_n767_;
  assign po115 = new_n768_;
  assign new_n842_ = ~new_n768_;
  assign po116 = new_n769_;
  assign new_n844_ = ~new_n769_;
  assign po117 = new_n770_;
  assign new_n846_ = ~new_n770_;
  assign new_n847_ = new_n771_;
  assign new_n848_ = new_n771_;
  assign new_n849_ = ~new_n772_;
  assign new_n850_ = pi029 & new_n751_ & new_n735_;
  assign new_n851_ = new_n722_ & pi027 & new_n433_ & pi191;
  assign new_n852_ = new_n660_ | new_n773_;
  assign new_n853_ = new_n661_ | new_n774_;
  assign new_n854_ = new_n662_ | new_n778_;
  assign new_n855_ = new_n663_ | new_n780_;
  assign new_n856_ = new_n664_ | new_n776_;
  assign new_n857_ = new_n665_ | new_n775_;
  assign new_n858_ = new_n666_ | new_n779_;
  assign new_n859_ = new_n667_ | new_n777_;
  assign new_n860_ = new_n668_ | new_n784_;
  assign new_n861_ = new_n669_ | new_n781_;
  assign new_n862_ = new_n670_ | new_n782_;
  assign new_n863_ = new_n671_ | new_n783_;
  assign new_n864_ = new_n672_ | new_n788_;
  assign new_n865_ = new_n673_ | new_n786_;
  assign new_n866_ = new_n675_ | new_n785_;
  assign new_n867_ = new_n676_ | new_n787_;
  assign new_n868_ = new_n677_ | new_n789_;
  assign new_n869_ = new_n802_ & new_n678_ & new_n729_;
  assign new_n870_ = new_n806_ & new_n679_ & new_n734_;
  assign new_n871_ = ~new_n794_ | ~new_n717_;
  assign new_n872_ = ~new_n796_ & ~new_n718_;
  assign new_n873_ = ~new_n795_ & ~new_n721_;
  assign new_n874_ = new_n800_ | new_n798_;
  assign new_n875_ = ~new_n723_ | ~new_n823_;
  assign new_n876_ = new_n801_ | new_n822_;
  assign new_n877_ = ~new_n852_ | ~new_n570_;
  assign new_n878_ = ~new_n853_ | ~new_n572_;
  assign new_n879_ = ~new_n857_ | ~new_n574_;
  assign new_n880_ = new_n803_ & new_n715_ & new_n689_;
  assign new_n881_ = ~new_n854_ | ~new_n576_;
  assign new_n882_ = ~new_n858_ | ~new_n578_;
  assign new_n883_ = ~new_n855_ | ~new_n579_;
  assign new_n884_ = ~new_n805_ | ~new_n804_;
  assign new_n885_ = ~new_n859_ | ~new_n581_;
  assign new_n886_ = ~new_n860_ | ~new_n583_;
  assign new_n887_ = ~new_n866_ | ~new_n585_;
  assign new_n888_ = ~new_n861_ | ~new_n587_;
  assign new_n889_ = ~new_n862_ | ~new_n589_;
  assign new_n890_ = ~new_n863_ | ~new_n591_;
  assign new_n891_ = new_n807_ & new_n716_ & new_n693_;
  assign new_n892_ = ~new_n867_ | ~new_n593_;
  assign new_n893_ = ~new_n864_ | ~new_n595_;
  assign new_n894_ = ~new_n868_ | ~new_n596_;
  assign new_n895_ = ~new_n865_ | ~new_n598_;
  assign new_n896_ = new_n738_ | new_n811_;
  assign new_n897_ = new_n810_ | new_n739_;
  assign new_n898_ = new_n813_ & pi198;
  assign new_n899_ = new_n813_ & new_n432_;
  assign new_n900_ = ~new_n813_;
  assign new_n901_ = new_n813_;
  assign po110 = ~new_n814_;
  assign new_n903_ = ~new_n696_ | ~new_n824_;
  assign new_n904_ = ~new_n744_ | ~new_n817_;
  assign new_n905_ = ~new_n746_ | ~new_n816_;
  assign new_n906_ = ~new_n747_ | ~new_n819_;
  assign new_n907_ = ~new_n749_ | ~new_n818_;
  assign new_n908_ = ~new_n752_ | ~new_n821_;
  assign new_n909_ = ~new_n754_ | ~new_n820_;
  assign new_n910_ = ~new_n755_ | ~new_n799_;
  assign new_n911_ = ~new_n825_;
  assign new_n912_ = ~new_n826_;
  assign new_n913_ = ~new_n827_;
  assign new_n914_ = ~new_n828_;
  assign new_n915_ = ~new_n829_;
  assign new_n916_ = ~new_n830_;
  assign new_n917_ = ~new_n831_;
  assign new_n918_ = ~new_n832_;
  assign new_n919_ = ~new_n832_ | ~new_n849_;
  assign new_n920_ = new_n834_;
  assign new_n921_ = new_n834_;
  assign new_n922_ = new_n834_;
  assign new_n923_ = new_n834_;
  assign new_n924_ = new_n836_;
  assign new_n925_ = new_n836_;
  assign new_n926_ = new_n836_;
  assign new_n927_ = ~new_n838_;
  assign new_n928_ = new_n840_;
  assign new_n929_ = new_n840_;
  assign new_n930_ = new_n842_;
  assign new_n931_ = new_n842_;
  assign new_n932_ = new_n844_;
  assign new_n933_ = new_n844_;
  assign new_n934_ = new_n846_;
  assign new_n935_ = new_n846_;
  assign new_n936_ = ~new_n847_;
  assign new_n937_ = ~new_n848_;
  assign new_n938_ = new_n808_ & pi029 & new_n751_;
  assign new_n939_ = new_n850_;
  assign new_n940_ = ~new_n850_;
  assign new_n941_ = ~new_n850_;
  assign new_n942_ = new_n850_;
  assign new_n943_ = ~new_n850_;
  assign po109 = ~new_n851_;
  assign new_n945_ = ~new_n852_;
  assign new_n946_ = ~new_n853_;
  assign new_n947_ = ~new_n854_;
  assign new_n948_ = ~new_n855_;
  assign new_n949_ = ~new_n857_;
  assign new_n950_ = ~new_n858_;
  assign new_n951_ = ~new_n859_;
  assign new_n952_ = ~new_n860_;
  assign new_n953_ = ~new_n861_;
  assign new_n954_ = ~new_n862_;
  assign new_n955_ = ~new_n863_;
  assign new_n956_ = ~new_n864_;
  assign new_n957_ = ~new_n865_;
  assign new_n958_ = ~new_n866_;
  assign new_n959_ = ~new_n867_;
  assign new_n960_ = ~new_n868_;
  assign new_n961_ = ~new_n880_ & ~new_n790_;
  assign new_n962_ = ~new_n869_ & ~new_n791_;
  assign new_n963_ = ~new_n891_ & ~new_n792_;
  assign new_n964_ = ~new_n870_ & ~new_n793_;
  assign new_n965_ = ~new_n871_;
  assign new_n966_ = ~new_n872_ | ~new_n873_;
  assign new_n967_ = ~new_n874_;
  assign new_n968_ = ~new_n910_ | ~new_n875_;
  assign new_n969_ = ~new_n876_;
  assign new_n970_ = ~new_n482_ | ~new_n945_;
  assign new_n971_ = ~new_n484_ | ~new_n946_;
  assign new_n972_ = ~new_n486_ | ~new_n949_;
  assign new_n973_ = ~new_n488_ | ~new_n947_;
  assign new_n974_ = ~new_n491_ | ~new_n950_;
  assign new_n975_ = ~new_n493_ | ~new_n948_;
  assign new_n976_ = ~new_n884_;
  assign new_n977_ = ~new_n495_ | ~new_n951_;
  assign new_n978_ = ~new_n497_ | ~new_n952_;
  assign new_n979_ = ~new_n499_ | ~new_n958_;
  assign new_n980_ = ~new_n501_ | ~new_n953_;
  assign new_n981_ = ~new_n503_ | ~new_n954_;
  assign new_n982_ = ~new_n505_ | ~new_n955_;
  assign new_n983_ = ~new_n507_ | ~new_n959_;
  assign new_n984_ = ~new_n509_ | ~new_n956_;
  assign new_n985_ = ~new_n511_ | ~new_n960_;
  assign new_n986_ = ~new_n513_ | ~new_n957_;
  assign new_n987_ = new_n737_ | new_n898_;
  assign po118 = new_n896_;
  assign po119 = new_n896_;
  assign po120 = new_n897_;
  assign po121 = new_n897_;
  assign po122 = new_n899_ | new_n741_;
  assign new_n993_ = ~new_n900_;
  assign new_n994_ = ~new_n901_;
  assign new_n995_ = ~new_n903_ | ~new_n815_;
  assign new_n996_ = new_n697_ & new_n941_;
  assign new_n997_ = new_n697_ & new_n940_;
  assign new_n998_ = ~new_n904_ | ~new_n905_;
  assign new_n999_ = new_n745_ & new_n941_;
  assign new_n1000_ = new_n745_ & new_n940_;
  assign new_n1001_ = ~new_n906_ | ~new_n907_;
  assign new_n1002_ = ~new_n908_ | ~new_n909_;
  assign new_n1003_ = new_n704_ & new_n941_;
  assign new_n1004_ = new_n704_ & new_n940_;
  assign new_n1005_ = ~new_n826_ | ~new_n936_;
  assign new_n1006_ = ~new_n827_ | ~new_n937_;
  assign new_n1007_ = ~new_n921_ | ~new_n915_;
  assign new_n1008_ = ~new_n923_ | ~new_n917_;
  assign new_n1009_ = ~new_n920_;
  assign new_n1010_ = ~new_n921_;
  assign new_n1011_ = ~new_n922_;
  assign new_n1012_ = ~new_n923_;
  assign new_n1013_ = ~new_n924_;
  assign new_n1014_ = ~new_n925_;
  assign new_n1015_ = ~new_n926_ | ~new_n927_;
  assign new_n1016_ = ~new_n926_;
  assign new_n1017_ = new_n765_ & new_n942_;
  assign new_n1018_ = new_n765_ & new_n939_;
  assign new_n1019_ = new_n767_ & new_n942_;
  assign new_n1020_ = new_n767_ & new_n939_;
  assign new_n1021_ = ~new_n928_;
  assign new_n1022_ = ~new_n929_;
  assign new_n1023_ = ~new_n930_;
  assign new_n1024_ = ~new_n931_;
  assign new_n1025_ = ~new_n932_;
  assign new_n1026_ = ~new_n933_;
  assign new_n1027_ = new_n770_ & new_n941_;
  assign new_n1028_ = new_n770_ & new_n940_;
  assign new_n1029_ = ~new_n934_;
  assign new_n1030_ = ~new_n935_;
  assign new_n1031_ = ~new_n847_ | ~new_n912_;
  assign new_n1032_ = ~new_n848_ | ~new_n913_;
  assign new_n1033_ = ~new_n772_ | ~new_n918_;
  assign new_n1034_ = new_n938_;
  assign new_n1035_ = new_n938_;
  assign new_n1036_ = ~new_n939_;
  assign new_n1037_ = ~new_n942_;
  assign new_n1038_ = new_n943_;
  assign new_n1039_ = new_n943_;
  assign new_n1040_ = ~new_n962_ | ~new_n961_;
  assign new_n1041_ = ~new_n964_ | ~new_n963_;
  assign new_n1042_ = ~new_n966_ | ~new_n965_;
  assign new_n1043_ = ~new_n966_;
  assign new_n1044_ = new_n874_ & new_n967_;
  assign new_n1045_ = ~new_n968_;
  assign new_n1046_ = new_n876_ & new_n969_;
  assign new_n1047_ = ~new_n877_ | ~new_n970_;
  assign new_n1048_ = ~new_n878_ | ~new_n971_;
  assign new_n1049_ = ~new_n879_ | ~new_n972_;
  assign new_n1050_ = ~new_n881_ | ~new_n973_;
  assign new_n1051_ = ~new_n882_ | ~new_n974_;
  assign new_n1052_ = ~new_n883_ | ~new_n975_;
  assign new_n1053_ = ~new_n885_ | ~new_n977_;
  assign new_n1054_ = ~new_n886_ | ~new_n978_;
  assign new_n1055_ = ~new_n887_ | ~new_n979_;
  assign new_n1056_ = ~new_n888_ | ~new_n980_;
  assign new_n1057_ = ~new_n889_ | ~new_n981_;
  assign new_n1058_ = ~new_n890_ | ~new_n982_;
  assign new_n1059_ = ~new_n892_ | ~new_n983_;
  assign new_n1060_ = ~new_n893_ | ~new_n984_;
  assign new_n1061_ = ~new_n894_ | ~new_n985_;
  assign new_n1062_ = ~new_n895_ | ~new_n986_;
  assign po123 = new_n987_;
  assign po124 = new_n987_;
  assign new_n1065_ = ~new_n995_;
  assign new_n1066_ = ~new_n998_;
  assign new_n1067_ = new_n1001_;
  assign new_n1068_ = new_n1001_;
  assign new_n1069_ = ~new_n1002_;
  assign new_n1070_ = ~new_n1005_ | ~new_n1031_;
  assign new_n1071_ = ~new_n1006_ | ~new_n1032_;
  assign new_n1072_ = ~new_n829_ | ~new_n1010_;
  assign new_n1073_ = ~new_n831_ | ~new_n1012_;
  assign new_n1074_ = ~new_n1033_ | ~new_n919_;
  assign new_n1075_ = new_n765_ & new_n1037_;
  assign new_n1076_ = new_n765_ & new_n1036_;
  assign new_n1077_ = ~new_n838_ | ~new_n1016_;
  assign new_n1078_ = new_n767_ & new_n1037_;
  assign new_n1079_ = new_n767_ & new_n1036_;
  assign new_n1080_ = ~new_n928_ | ~new_n1023_;
  assign new_n1081_ = ~new_n929_ | ~new_n1024_;
  assign new_n1082_ = new_n768_ & new_n1037_;
  assign new_n1083_ = new_n768_ & new_n1036_;
  assign new_n1084_ = ~new_n930_ | ~new_n1021_;
  assign new_n1085_ = ~new_n931_ | ~new_n1022_;
  assign new_n1086_ = new_n769_ & new_n1037_;
  assign new_n1087_ = new_n769_ & new_n1036_;
  assign new_n1088_ = ~new_n932_ | ~new_n1029_;
  assign new_n1089_ = ~new_n933_ | ~new_n1030_;
  assign new_n1090_ = ~new_n934_ | ~new_n1025_;
  assign new_n1091_ = ~new_n935_ | ~new_n1026_;
  assign new_n1092_ = new_n1034_;
  assign new_n1093_ = new_n1034_;
  assign new_n1094_ = new_n1035_;
  assign new_n1095_ = new_n1035_;
  assign new_n1096_ = new_n1038_;
  assign new_n1097_ = new_n1038_;
  assign new_n1098_ = new_n1038_;
  assign new_n1099_ = new_n1039_;
  assign new_n1100_ = new_n1039_;
  assign new_n1101_ = new_n1039_;
  assign new_n1102_ = ~new_n1040_;
  assign new_n1103_ = ~new_n1041_;
  assign new_n1104_ = ~new_n871_ | ~new_n1043_;
  assign new_n1105_ = new_n1044_ | new_n967_;
  assign new_n1106_ = ~new_n968_ | ~new_n1069_;
  assign new_n1107_ = ~new_n1040_ | ~new_n725_;
  assign new_n1108_ = new_n1046_ | new_n969_;
  assign new_n1109_ = ~new_n1047_;
  assign new_n1110_ = ~new_n1048_;
  assign new_n1111_ = ~new_n1049_;
  assign new_n1112_ = ~new_n1050_;
  assign new_n1113_ = new_n401_ & new_n1097_;
  assign new_n1114_ = new_n401_ & new_n1100_;
  assign new_n1115_ = ~new_n1051_;
  assign new_n1116_ = new_n406_ & new_n1097_;
  assign new_n1117_ = new_n406_ & new_n1100_;
  assign new_n1118_ = ~new_n1052_;
  assign new_n1119_ = ~new_n1041_ | ~new_n976_;
  assign new_n1120_ = new_n408_ & new_n1097_;
  assign new_n1121_ = new_n408_ & new_n1100_;
  assign new_n1122_ = ~new_n1053_;
  assign new_n1123_ = new_n410_ & new_n1097_;
  assign new_n1124_ = new_n410_ & new_n1100_;
  assign new_n1125_ = ~new_n1054_;
  assign new_n1126_ = new_n412_ & new_n1096_;
  assign new_n1127_ = new_n412_ & new_n1099_;
  assign new_n1128_ = ~new_n1055_;
  assign new_n1129_ = new_n414_ & new_n1096_;
  assign new_n1130_ = new_n414_ & new_n1099_;
  assign new_n1131_ = ~new_n1056_;
  assign new_n1132_ = new_n416_ & new_n1096_;
  assign new_n1133_ = new_n416_ & new_n1099_;
  assign new_n1134_ = ~new_n1057_;
  assign new_n1135_ = new_n418_ & new_n1096_;
  assign new_n1136_ = new_n418_ & new_n1099_;
  assign new_n1137_ = ~new_n1058_;
  assign new_n1138_ = new_n420_ & new_n1098_;
  assign new_n1139_ = new_n420_ & new_n1101_;
  assign new_n1140_ = ~new_n1059_;
  assign new_n1141_ = new_n422_ & new_n1098_;
  assign new_n1142_ = new_n422_ & new_n1101_;
  assign new_n1143_ = ~new_n1060_;
  assign new_n1144_ = new_n425_ & new_n1101_;
  assign new_n1145_ = new_n425_ & new_n1098_;
  assign new_n1146_ = ~new_n1061_;
  assign new_n1147_ = new_n427_ & new_n1098_;
  assign new_n1148_ = new_n427_ & new_n1101_;
  assign new_n1149_ = ~new_n1062_;
  assign new_n1150_ = ~new_n1074_ | ~new_n993_;
  assign new_n1151_ = new_n1068_ & new_n998_ & new_n995_;
  assign new_n1152_ = new_n1067_ & new_n1066_ & new_n1065_;
  assign new_n1153_ = new_n996_ & new_n1092_;
  assign new_n1154_ = new_n997_ & new_n1093_;
  assign new_n1155_ = new_n999_ & new_n1092_;
  assign new_n1156_ = new_n1000_ & new_n1093_;
  assign new_n1157_ = ~new_n1067_;
  assign new_n1158_ = ~new_n1068_;
  assign new_n1159_ = ~new_n1002_ | ~new_n1045_;
  assign new_n1160_ = new_n1003_ & new_n1092_;
  assign new_n1161_ = new_n1004_ & new_n1093_;
  assign new_n1162_ = ~new_n1070_;
  assign new_n1163_ = ~new_n1071_;
  assign new_n1164_ = ~new_n1072_ | ~new_n1007_;
  assign new_n1165_ = ~new_n1073_ | ~new_n1008_;
  assign new_n1166_ = ~new_n1074_;
  assign new_n1167_ = ~new_n1015_ | ~new_n1077_;
  assign new_n1168_ = new_n1075_ | new_n1017_;
  assign new_n1169_ = new_n1076_ | new_n1018_;
  assign new_n1170_ = new_n1078_ | new_n1019_;
  assign new_n1171_ = new_n1079_ | new_n1020_;
  assign new_n1172_ = ~new_n1080_ | ~new_n1084_;
  assign new_n1173_ = ~new_n1081_ | ~new_n1085_;
  assign new_n1174_ = ~new_n1088_ | ~new_n1090_;
  assign new_n1175_ = ~new_n1089_ | ~new_n1091_;
  assign new_n1176_ = new_n1027_ & new_n1092_;
  assign new_n1177_ = new_n1028_ & new_n1093_;
  assign new_n1178_ = ~new_n1096_;
  assign new_n1179_ = ~new_n1098_;
  assign new_n1180_ = ~new_n1099_;
  assign new_n1181_ = ~new_n1101_;
  assign new_n1182_ = new_n1082_ & new_n552_;
  assign new_n1183_ = new_n1086_ & new_n552_;
  assign new_n1184_ = new_n1083_ & new_n553_;
  assign new_n1185_ = new_n1087_ & new_n553_;
  assign new_n1186_ = ~new_n1104_ | ~new_n1042_;
  assign po125 = ~new_n1105_ | ~new_n1108_;
  assign new_n1188_ = ~new_n1159_ | ~new_n1106_;
  assign new_n1189_ = ~new_n687_ | ~new_n1102_;
  assign new_n1190_ = new_n392_ & new_n1178_;
  assign new_n1191_ = new_n392_ & new_n1180_;
  assign new_n1192_ = new_n394_ & new_n1178_;
  assign new_n1193_ = new_n394_ & new_n1180_;
  assign new_n1194_ = new_n1118_ & new_n1115_ & new_n1112_ & new_n1110_ & new_n1111_;
  assign new_n1195_ = new_n396_ & new_n1179_;
  assign new_n1196_ = new_n396_ & new_n1181_;
  assign new_n1197_ = new_n398_ & new_n1179_;
  assign new_n1198_ = new_n398_ & new_n1181_;
  assign new_n1199_ = new_n401_ & new_n1179_;
  assign new_n1200_ = new_n401_ & new_n1181_;
  assign new_n1201_ = new_n406_ & new_n1179_;
  assign new_n1202_ = new_n406_ & new_n1181_;
  assign new_n1203_ = ~new_n884_ | ~new_n1103_;
  assign new_n1204_ = new_n1134_ & new_n1131_ & new_n1128_ & new_n1122_ & new_n1125_;
  assign new_n1205_ = new_n1149_ & new_n1146_ & new_n1143_ & new_n1137_ & new_n1140_;
  assign new_n1206_ = ~new_n900_ | ~new_n1166_;
  assign new_n1207_ = new_n1157_ & new_n995_ & new_n1066_;
  assign new_n1208_ = ~new_n1153_;
  assign new_n1209_ = ~new_n1154_;
  assign new_n1210_ = new_n1158_ & new_n1065_ & new_n998_;
  assign new_n1211_ = ~new_n1155_;
  assign new_n1212_ = ~new_n1156_;
  assign new_n1213_ = ~new_n1160_;
  assign new_n1214_ = ~new_n1161_;
  assign new_n1215_ = ~new_n1164_;
  assign new_n1216_ = new_n1165_;
  assign new_n1217_ = new_n1165_;
  assign new_n1218_ = new_n1167_;
  assign new_n1219_ = new_n1167_;
  assign new_n1220_ = ~new_n1172_;
  assign new_n1221_ = ~new_n1173_;
  assign new_n1222_ = ~new_n1174_;
  assign new_n1223_ = ~new_n1175_;
  assign new_n1224_ = ~new_n1176_;
  assign new_n1225_ = ~new_n1177_;
  assign new_n1226_ = new_n1116_ & new_n1094_;
  assign new_n1227_ = new_n1120_ & new_n1094_;
  assign new_n1228_ = new_n1123_ & new_n1094_;
  assign new_n1229_ = new_n1113_ & new_n1094_;
  assign new_n1230_ = new_n1117_ & new_n1095_;
  assign new_n1231_ = new_n1121_ & new_n1095_;
  assign new_n1232_ = new_n1124_ & new_n1095_;
  assign new_n1233_ = new_n1114_ & new_n1095_;
  assign new_n1234_ = new_n856_ & new_n1109_;
  assign new_n1235_ = new_n1126_ & new_n550_;
  assign new_n1236_ = new_n1129_ & new_n550_;
  assign new_n1237_ = new_n1127_ & new_n551_;
  assign new_n1238_ = new_n1130_ & new_n551_;
  assign new_n1239_ = new_n1168_ & new_n552_;
  assign new_n1240_ = new_n1170_ & new_n552_;
  assign new_n1241_ = ~new_n1182_;
  assign new_n1242_ = ~new_n1183_;
  assign new_n1243_ = new_n1169_ & new_n553_;
  assign new_n1244_ = new_n1171_ & new_n553_;
  assign new_n1245_ = ~new_n1184_;
  assign new_n1246_ = ~new_n1185_;
  assign new_n1247_ = ~new_n1186_;
  assign new_n1248_ = ~new_n1188_;
  assign new_n1249_ = ~new_n1189_ | ~new_n1107_;
  assign new_n1250_ = new_n1234_ & new_n1194_;
  assign new_n1251_ = ~new_n1203_ | ~new_n1119_;
  assign new_n1252_ = new_n1204_ & new_n1205_;
  assign new_n1253_ = new_n1190_ | new_n1132_;
  assign new_n1254_ = new_n1191_ | new_n1133_;
  assign new_n1255_ = new_n1192_ | new_n1135_;
  assign new_n1256_ = new_n1193_ | new_n1136_;
  assign new_n1257_ = new_n1195_ | new_n1138_;
  assign new_n1258_ = new_n1196_ | new_n1139_;
  assign new_n1259_ = new_n1197_ | new_n1141_;
  assign new_n1260_ = new_n1198_ | new_n1142_;
  assign new_n1261_ = new_n1200_ | new_n1144_;
  assign new_n1262_ = new_n1199_ | new_n1145_;
  assign new_n1263_ = new_n1201_ | new_n1147_;
  assign new_n1264_ = new_n1202_ | new_n1148_;
  assign new_n1265_ = ~new_n1150_ | ~new_n1206_;
  assign new_n1266_ = new_n1216_ & new_n1071_ & new_n901_;
  assign new_n1267_ = new_n1217_ & new_n1163_ & new_n994_;
  assign new_n1268_ = ~new_n1210_ & ~new_n1151_;
  assign new_n1269_ = ~new_n1207_ & ~new_n1152_;
  assign new_n1270_ = new_n1226_ & new_n1208_;
  assign new_n1271_ = new_n1208_;
  assign new_n1272_ = new_n1230_ & new_n1209_;
  assign new_n1273_ = new_n1209_;
  assign new_n1274_ = new_n1229_ & new_n1211_;
  assign new_n1275_ = new_n1211_;
  assign new_n1276_ = new_n1233_ & new_n1212_;
  assign new_n1277_ = new_n1212_;
  assign new_n1278_ = new_n1227_ & new_n1213_;
  assign new_n1279_ = new_n1213_;
  assign new_n1280_ = new_n1231_ & new_n1214_;
  assign new_n1281_ = new_n1214_;
  assign new_n1282_ = new_n1219_ & new_n1164_ & new_n1070_;
  assign new_n1283_ = new_n1218_ & new_n1215_ & new_n1162_;
  assign new_n1284_ = ~new_n1216_;
  assign new_n1285_ = ~new_n1217_;
  assign new_n1286_ = ~new_n1218_;
  assign new_n1287_ = ~new_n1219_;
  assign new_n1288_ = ~new_n1172_ | ~new_n1222_;
  assign new_n1289_ = ~new_n1173_ | ~new_n1223_;
  assign new_n1290_ = ~new_n1174_ | ~new_n1220_;
  assign new_n1291_ = ~new_n1175_ | ~new_n1221_;
  assign new_n1292_ = new_n1224_ & new_n1228_;
  assign new_n1293_ = new_n1224_;
  assign new_n1294_ = new_n1225_ & new_n1232_;
  assign new_n1295_ = new_n1225_;
  assign new_n1296_ = new_n1226_;
  assign new_n1297_ = new_n1227_;
  assign new_n1298_ = new_n1228_;
  assign new_n1299_ = new_n1229_;
  assign new_n1300_ = new_n1230_;
  assign new_n1301_ = new_n1231_;
  assign new_n1302_ = new_n1232_;
  assign new_n1303_ = new_n1233_;
  assign new_n1304_ = new_n1235_ & new_n1242_;
  assign new_n1305_ = new_n1235_;
  assign new_n1306_ = new_n1236_ & new_n1241_;
  assign new_n1307_ = new_n1236_;
  assign new_n1308_ = new_n1237_ & new_n1246_;
  assign new_n1309_ = new_n1237_;
  assign new_n1310_ = new_n1238_ & new_n1245_;
  assign new_n1311_ = new_n1238_;
  assign new_n1312_ = ~new_n1239_;
  assign new_n1313_ = ~new_n1240_;
  assign new_n1314_ = new_n1241_;
  assign new_n1315_ = new_n1242_;
  assign new_n1316_ = ~new_n1243_;
  assign new_n1317_ = ~new_n1244_;
  assign new_n1318_ = new_n1245_;
  assign new_n1319_ = new_n1246_;
  assign po127 = ~new_n1249_;
  assign po128 = ~new_n1251_;
  assign new_n1322_ = new_n1257_;
  assign new_n1323_ = new_n1258_;
  assign new_n1324_ = new_n1259_;
  assign new_n1325_ = new_n1260_;
  assign new_n1326_ = new_n1261_;
  assign new_n1327_ = new_n1262_;
  assign new_n1328_ = ~new_n1265_;
  assign new_n1329_ = new_n1285_ & new_n901_ & new_n1163_;
  assign new_n1330_ = new_n1284_ & new_n994_ & new_n1071_;
  assign new_n1331_ = ~new_n1269_ | ~new_n1268_;
  assign new_n1332_ = ~new_n1271_;
  assign new_n1333_ = ~new_n1273_;
  assign new_n1334_ = ~new_n1275_;
  assign new_n1335_ = ~new_n1277_;
  assign new_n1336_ = ~new_n1279_;
  assign new_n1337_ = ~new_n1281_;
  assign new_n1338_ = ~new_n1265_ | ~new_n911_;
  assign new_n1339_ = new_n1286_ & new_n1070_ & new_n1215_;
  assign new_n1340_ = new_n1287_ & new_n1162_ & new_n1164_;
  assign new_n1341_ = new_n1262_ & new_n759_;
  assign new_n1342_ = new_n1261_ & new_n759_;
  assign new_n1343_ = new_n1259_ & new_n834_;
  assign new_n1344_ = new_n1260_ & new_n834_;
  assign new_n1345_ = new_n1257_ & new_n836_;
  assign new_n1346_ = new_n1258_ & new_n836_;
  assign new_n1347_ = ~new_n1288_ | ~new_n1290_;
  assign new_n1348_ = ~new_n1289_ | ~new_n1291_;
  assign new_n1349_ = ~new_n1293_;
  assign new_n1350_ = ~new_n1295_;
  assign new_n1351_ = new_n1263_ & new_n771_;
  assign new_n1352_ = new_n1264_ & new_n771_;
  assign new_n1353_ = ~new_n1296_;
  assign new_n1354_ = ~new_n1297_;
  assign new_n1355_ = ~new_n1298_;
  assign new_n1356_ = ~new_n1299_;
  assign new_n1357_ = ~new_n1300_;
  assign new_n1358_ = ~new_n1301_;
  assign new_n1359_ = ~new_n1302_;
  assign new_n1360_ = ~new_n1303_;
  assign new_n1361_ = new_n1247_ & pi009;
  assign new_n1362_ = new_n674_ & new_n1252_ & new_n1250_;
  assign new_n1363_ = ~new_n1305_;
  assign new_n1364_ = ~new_n1307_;
  assign new_n1365_ = new_n1253_ & new_n550_;
  assign new_n1366_ = new_n1255_ & new_n550_;
  assign new_n1367_ = ~new_n1309_;
  assign new_n1368_ = ~new_n1311_;
  assign new_n1369_ = new_n1254_ & new_n551_;
  assign new_n1370_ = new_n1256_ & new_n551_;
  assign new_n1371_ = new_n1312_;
  assign new_n1372_ = new_n1313_;
  assign new_n1373_ = ~new_n1314_;
  assign new_n1374_ = ~new_n1315_;
  assign new_n1375_ = new_n1316_;
  assign new_n1376_ = new_n1317_;
  assign new_n1377_ = ~new_n1318_;
  assign new_n1378_ = ~new_n1319_;
  assign new_n1379_ = ~new_n1331_ | ~new_n1248_;
  assign new_n1380_ = ~new_n1322_;
  assign new_n1381_ = ~new_n1323_;
  assign new_n1382_ = ~new_n1324_;
  assign new_n1383_ = ~new_n1325_;
  assign new_n1384_ = ~new_n1326_;
  assign new_n1385_ = ~new_n1327_;
  assign new_n1386_ = ~new_n1330_ & ~new_n1266_;
  assign new_n1387_ = ~new_n1329_ & ~new_n1267_;
  assign new_n1388_ = ~new_n1331_;
  assign new_n1389_ = ~new_n1271_ | ~new_n1353_;
  assign new_n1390_ = ~new_n1273_ | ~new_n1357_;
  assign new_n1391_ = ~new_n1275_ | ~new_n1356_;
  assign new_n1392_ = ~new_n1277_ | ~new_n1360_;
  assign new_n1393_ = ~new_n1279_ | ~new_n1354_;
  assign new_n1394_ = ~new_n1281_ | ~new_n1358_;
  assign new_n1395_ = ~new_n825_ | ~new_n1328_;
  assign new_n1396_ = ~new_n1340_ & ~new_n1282_;
  assign new_n1397_ = ~new_n1339_ & ~new_n1283_;
  assign new_n1398_ = ~new_n1326_ | ~new_n914_;
  assign new_n1399_ = ~new_n1327_ | ~new_n916_;
  assign new_n1400_ = ~new_n1325_ | ~new_n1009_;
  assign new_n1401_ = ~new_n1324_ | ~new_n1011_;
  assign new_n1402_ = ~new_n1323_ | ~new_n1013_;
  assign new_n1403_ = ~new_n1322_ | ~new_n1014_;
  assign new_n1404_ = ~new_n1347_;
  assign new_n1405_ = ~new_n1348_;
  assign new_n1406_ = ~new_n1293_ | ~new_n1355_;
  assign new_n1407_ = ~new_n1295_ | ~new_n1359_;
  assign new_n1408_ = ~new_n1296_ | ~new_n1332_;
  assign new_n1409_ = ~new_n1297_ | ~new_n1336_;
  assign new_n1410_ = ~new_n1298_ | ~new_n1349_;
  assign new_n1411_ = ~new_n1299_ | ~new_n1334_;
  assign new_n1412_ = ~new_n1300_ | ~new_n1333_;
  assign new_n1413_ = ~new_n1301_ | ~new_n1337_;
  assign new_n1414_ = ~new_n1302_ | ~new_n1350_;
  assign new_n1415_ = ~new_n1303_ | ~new_n1335_;
  assign new_n1416_ = ~new_n1361_;
  assign po126 = new_n1361_;
  assign po130 = ~new_n1362_;
  assign po129 = new_n1362_;
  assign new_n1420_ = ~new_n1305_ | ~new_n1374_;
  assign new_n1421_ = ~new_n1307_ | ~new_n1373_;
  assign new_n1422_ = new_n1365_;
  assign new_n1423_ = new_n1366_;
  assign new_n1424_ = ~new_n1309_ | ~new_n1378_;
  assign new_n1425_ = ~new_n1311_ | ~new_n1377_;
  assign new_n1426_ = new_n1369_;
  assign new_n1427_ = new_n1370_;
  assign new_n1428_ = ~new_n1371_;
  assign new_n1429_ = new_n1366_ & new_n1312_;
  assign new_n1430_ = new_n1365_ & new_n1313_;
  assign new_n1431_ = ~new_n1372_;
  assign new_n1432_ = ~new_n1314_ | ~new_n1364_;
  assign new_n1433_ = ~new_n1315_ | ~new_n1363_;
  assign new_n1434_ = ~new_n1375_;
  assign new_n1435_ = new_n1370_ & new_n1316_;
  assign new_n1436_ = new_n1369_ & new_n1317_;
  assign new_n1437_ = ~new_n1376_;
  assign new_n1438_ = ~new_n1318_ | ~new_n1368_;
  assign new_n1439_ = ~new_n1319_ | ~new_n1367_;
  assign new_n1440_ = ~new_n1188_ | ~new_n1388_;
  assign new_n1441_ = ~new_n1387_ | ~new_n1386_;
  assign new_n1442_ = ~new_n1389_ | ~new_n1408_;
  assign new_n1443_ = ~new_n1390_ | ~new_n1412_;
  assign new_n1444_ = ~new_n1391_ | ~new_n1411_;
  assign new_n1445_ = ~new_n1392_ | ~new_n1415_;
  assign new_n1446_ = ~new_n1393_ | ~new_n1409_;
  assign new_n1447_ = ~new_n1394_ | ~new_n1413_;
  assign new_n1448_ = ~new_n1338_ | ~new_n1395_;
  assign new_n1449_ = ~new_n1397_ | ~new_n1396_;
  assign new_n1450_ = ~new_n828_ | ~new_n1384_;
  assign new_n1451_ = ~new_n830_ | ~new_n1385_;
  assign new_n1452_ = ~new_n920_ | ~new_n1383_;
  assign new_n1453_ = ~new_n922_ | ~new_n1382_;
  assign new_n1454_ = ~new_n924_ | ~new_n1381_;
  assign new_n1455_ = ~new_n925_ | ~new_n1380_;
  assign new_n1456_ = ~new_n1406_ | ~new_n1410_;
  assign new_n1457_ = ~new_n1407_ | ~new_n1414_;
  assign new_n1458_ = ~new_n1433_ | ~new_n1420_;
  assign new_n1459_ = ~new_n1432_ | ~new_n1421_;
  assign new_n1460_ = ~new_n1422_ | ~new_n1431_;
  assign new_n1461_ = ~new_n1422_;
  assign new_n1462_ = ~new_n1423_ | ~new_n1428_;
  assign new_n1463_ = ~new_n1423_;
  assign new_n1464_ = ~new_n1439_ | ~new_n1424_;
  assign new_n1465_ = ~new_n1438_ | ~new_n1425_;
  assign new_n1466_ = ~new_n1426_ | ~new_n1437_;
  assign new_n1467_ = ~new_n1426_;
  assign new_n1468_ = ~new_n1427_ | ~new_n1434_;
  assign new_n1469_ = ~new_n1427_;
  assign new_n1470_ = ~new_n1440_ | ~new_n1379_;
  assign new_n1471_ = new_n1448_ & new_n432_;
  assign new_n1472_ = ~new_n1441_;
  assign new_n1473_ = new_n1444_ & new_n1270_;
  assign new_n1474_ = new_n1444_ & new_n1446_ & new_n1442_ & new_n1456_;
  assign new_n1475_ = new_n1445_ & new_n1272_;
  assign new_n1476_ = new_n1445_ & new_n1447_ & new_n1443_ & new_n1457_;
  assign new_n1477_ = new_n1278_ & new_n1442_ & new_n1444_;
  assign new_n1478_ = new_n1280_ & new_n1443_ & new_n1445_;
  assign new_n1479_ = ~new_n1449_;
  assign new_n1480_ = ~new_n1450_ | ~new_n1398_;
  assign new_n1481_ = ~new_n1451_ | ~new_n1399_;
  assign new_n1482_ = ~new_n1452_ | ~new_n1400_;
  assign new_n1483_ = ~new_n1453_ | ~new_n1401_;
  assign new_n1484_ = ~new_n1454_ | ~new_n1402_;
  assign new_n1485_ = ~new_n1455_ | ~new_n1403_;
  assign new_n1486_ = ~new_n1449_ | ~new_n1404_;
  assign new_n1487_ = ~new_n1441_ | ~new_n1405_;
  assign new_n1488_ = new_n1442_ & new_n1292_ & new_n1446_ & new_n1444_;
  assign new_n1489_ = new_n1443_ & new_n1294_ & new_n1447_ & new_n1445_;
  assign new_n1490_ = new_n1458_ & new_n1306_;
  assign new_n1491_ = new_n1464_ & new_n1310_;
  assign new_n1492_ = ~new_n1371_ | ~new_n1463_;
  assign new_n1493_ = new_n1430_ & new_n1459_ & new_n1458_;
  assign new_n1494_ = ~new_n1372_ | ~new_n1461_;
  assign new_n1495_ = ~new_n1375_ | ~new_n1469_;
  assign new_n1496_ = new_n1436_ & new_n1465_ & new_n1464_;
  assign new_n1497_ = ~new_n1376_ | ~new_n1467_;
  assign new_n1498_ = ~new_n1470_;
  assign po131 = new_n1471_ | new_n742_;
  assign new_n1500_ = ~new_n1474_;
  assign new_n1501_ = ~new_n1476_;
  assign new_n1502_ = new_n1488_ | new_n1477_ | new_n1274_ | new_n1473_;
  assign new_n1503_ = new_n1489_ | new_n1478_ | new_n1276_ | new_n1475_;
  assign new_n1504_ = new_n1483_ & new_n1341_;
  assign new_n1505_ = new_n1482_ & new_n1342_;
  assign new_n1506_ = ~new_n1347_ | ~new_n1479_;
  assign new_n1507_ = ~new_n1348_ | ~new_n1472_;
  assign new_n1508_ = new_n1351_ & new_n1481_ & new_n1483_;
  assign new_n1509_ = new_n1352_ & new_n1480_ & new_n1482_;
  assign new_n1510_ = ~new_n1494_ | ~new_n1460_;
  assign new_n1511_ = ~new_n1492_ | ~new_n1462_;
  assign new_n1512_ = ~new_n1497_ | ~new_n1466_;
  assign new_n1513_ = ~new_n1495_ | ~new_n1468_;
  assign new_n1514_ = ~new_n1502_;
  assign new_n1515_ = ~new_n1503_;
  assign new_n1516_ = new_n1508_ | new_n1343_ | new_n1504_;
  assign new_n1517_ = new_n1509_ | new_n1344_ | new_n1505_;
  assign new_n1518_ = new_n1459_ & new_n1345_ & new_n1458_ & new_n1511_ & new_n1510_;
  assign new_n1519_ = new_n1465_ & new_n1346_ & new_n1464_ & new_n1513_ & new_n1512_;
  assign new_n1520_ = ~new_n1506_ | ~new_n1486_;
  assign new_n1521_ = ~new_n1507_ | ~new_n1487_;
  assign new_n1522_ = new_n1498_ & new_n544_;
  assign new_n1523_ = new_n1511_ & new_n1458_ & new_n1510_ & new_n1459_ & new_n1485_;
  assign new_n1524_ = new_n1513_ & new_n1464_ & new_n1512_ & new_n1465_ & new_n1484_;
  assign new_n1525_ = new_n1459_ & new_n1429_ & new_n1510_ & new_n1458_;
  assign new_n1526_ = new_n1465_ & new_n1435_ & new_n1512_ & new_n1464_;
  assign new_n1527_ = new_n1521_ & pi198;
  assign new_n1528_ = ~new_n1514_ | ~new_n1500_;
  assign new_n1529_ = ~new_n1515_ | ~new_n1501_;
  assign new_n1530_ = new_n1523_ & new_n1516_;
  assign new_n1531_ = new_n1524_ & new_n1517_;
  assign new_n1532_ = ~new_n1520_;
  assign po132 = new_n1522_;
  assign new_n1534_ = ~new_n1522_;
  assign new_n1535_ = new_n1518_ | new_n1525_ | new_n1493_ | new_n1304_ | new_n1490_;
  assign new_n1536_ = new_n1519_ | new_n1526_ | new_n1496_ | new_n1308_ | new_n1491_;
  assign new_n1537_ = new_n809_ | new_n1527_;
  assign new_n1538_ = new_n1535_ | new_n1530_;
  assign new_n1539_ = new_n1536_ | new_n1531_;
  assign new_n1540_ = new_n1532_ & new_n544_;
  assign po133 = new_n1537_;
  assign po134 = new_n1537_;
  assign new_n1543_ = new_n1528_ & new_n1538_;
  assign new_n1544_ = new_n1529_ & new_n1539_;
  assign new_n1545_ = ~new_n1538_;
  assign new_n1546_ = ~new_n1539_;
  assign po135 = new_n1540_;
  assign new_n1548_ = ~new_n1540_;
  assign new_n1549_ = new_n1249_ & new_n1534_ & new_n1548_;
  assign new_n1550_ = new_n1502_ & new_n1545_;
  assign new_n1551_ = new_n1503_ & new_n1546_;
  assign new_n1552_ = new_n1550_ | new_n1543_;
  assign new_n1553_ = new_n1551_ | new_n1544_;
  assign new_n1554_ = ~new_n1553_ | ~new_n1552_;
  assign po136 = new_n1553_;
  assign new_n1556_ = new_n1554_ & new_n1552_;
  assign new_n1557_ = new_n1553_ & new_n1554_;
  assign new_n1558_ = new_n1557_ | new_n1556_;
  assign new_n1559_ = ~new_n1558_;
  assign new_n1560_ = new_n1558_ & new_n1559_;
  assign new_n1561_ = new_n1560_ | new_n1559_;
  assign new_n1562_ = new_n1561_ & new_n1251_ & new_n1416_;
  assign po137 = ~new_n1561_;
  assign new_n1564_ = new_n722_ & new_n1549_ & new_n1562_;
  assign po139 = ~new_n1564_;
  assign po138 = new_n1564_;
  assign po000 = pi114;
  assign po001 = pi115;
  assign po002 = pi116;
  assign po003 = pi117;
  assign po004 = pi118;
  assign po005 = pi119;
  assign po006 = pi120;
  assign po007 = pi121;
  assign po008 = pi122;
  assign po009 = pi123;
  assign po010 = pi124;
  assign po011 = pi125;
  assign po012 = pi126;
  assign po013 = pi127;
  assign po014 = pi128;
  assign po015 = pi129;
  assign po016 = pi130;
  assign po017 = pi131;
  assign po018 = pi132;
  assign po019 = pi133;
  assign po020 = pi134;
  assign po021 = pi135;
  assign po022 = pi136;
  assign po023 = pi137;
  assign po024 = pi138;
  assign po025 = pi139;
  assign po026 = pi140;
  assign po027 = pi141;
  assign po028 = pi142;
  assign po029 = pi143;
  assign po030 = pi144;
  assign po031 = pi145;
  assign po032 = pi146;
  assign po033 = pi147;
  assign po034 = pi148;
  assign po035 = pi149;
  assign po036 = pi150;
  assign po037 = pi151;
  assign po038 = pi152;
  assign po039 = pi153;
  assign po040 = pi154;
  assign po041 = pi155;
  assign po042 = pi156;
  assign po043 = pi157;
  assign po044 = pi158;
  assign po045 = pi159;
  assign po046 = pi160;
  assign po047 = pi161;
  assign po048 = pi162;
  assign po049 = pi163;
  assign po050 = pi164;
  assign po051 = pi165;
  assign po052 = pi166;
  assign po053 = pi167;
  assign po054 = pi168;
  assign po055 = pi169;
  assign po056 = pi170;
  assign po057 = pi171;
  assign po058 = pi172;
  assign po059 = pi173;
  assign po060 = pi174;
  assign po061 = pi175;
  assign po062 = pi176;
  assign po063 = pi177;
  assign po064 = pi178;
  assign po065 = pi179;
  assign po066 = pi180;
  assign po067 = pi181;
  assign po068 = pi182;
  assign po069 = pi183;
  assign po070 = pi184;
  assign po071 = pi185;
  assign po072 = pi186;
  assign po073 = pi187;
  assign po074 = pi188;
  assign po075 = pi189;
endmodule


