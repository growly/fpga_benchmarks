// Benchmark "i4" written by ABC on Thu Mar 19 13:02:36 2020

module i4 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191,
    po0, po1, po2, po3, po4, po5  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191;
  output po0, po1, po2, po3, po4, po5;
  wire new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_;
  assign po0 = pi000 & pi001;
  assign po1 = pi002 & pi003;
  assign new_n201_ = pi004 & pi005;
  assign new_n202_ = pi006 & pi007;
  assign new_n203_ = pi008 & pi009;
  assign new_n204_ = pi010 & pi011;
  assign new_n205_ = pi012 & pi013;
  assign new_n206_ = pi014 & pi015;
  assign new_n207_ = pi016 & pi017;
  assign new_n208_ = pi018 & pi019;
  assign new_n209_ = pi020 & pi021;
  assign new_n210_ = pi022 & pi023;
  assign new_n211_ = pi024 & pi025;
  assign new_n212_ = pi026 & pi027;
  assign new_n213_ = pi028 & pi029;
  assign new_n214_ = pi030 & pi031;
  assign new_n215_ = pi032 & pi033;
  assign new_n216_ = pi034 & pi035;
  assign new_n217_ = pi038 & pi036 & pi037;
  assign new_n218_ = pi036 & pi041 & pi039 & pi040;
  assign new_n219_ = pi039 & pi044 & pi043 & pi042 & pi036;
  assign new_n220_ = pi047 & pi045 & pi046;
  assign new_n221_ = pi045 & pi050 & pi048 & pi049;
  assign new_n222_ = pi048 & pi053 & pi052 & pi051 & pi045;
  assign new_n223_ = pi056 & pi054 & pi055;
  assign new_n224_ = pi054 & pi059 & pi057 & pi058;
  assign new_n225_ = pi057 & pi062 & pi061 & pi060 & pi054;
  assign new_n226_ = pi065 & pi063 & pi064;
  assign new_n227_ = pi063 & pi068 & pi066 & pi067;
  assign new_n228_ = pi066 & pi071 & pi070 & pi069 & pi063;
  assign new_n229_ = new_n202_ | new_n221_ | new_n222_ | new_n220_;
  assign new_n230_ = new_n203_ | new_n224_ | new_n225_ | new_n223_;
  assign new_n231_ = new_n204_ | new_n227_ | new_n228_ | new_n226_;
  assign new_n232_ = pi074 & pi072 & pi073;
  assign new_n233_ = pi072 & pi077 & pi075 & pi076;
  assign new_n234_ = pi075 & pi080 & pi079 & pi078 & pi072;
  assign new_n235_ = pi083 & pi081 & pi082;
  assign new_n236_ = pi081 & pi086 & pi084 & pi085;
  assign new_n237_ = pi084 & pi089 & pi088 & pi087 & pi081;
  assign new_n238_ = pi092 & pi090 & pi091;
  assign new_n239_ = pi090 & pi095 & pi093 & pi094;
  assign new_n240_ = pi093 & pi098 & pi097 & pi096 & pi090;
  assign new_n241_ = pi101 & pi099 & pi100;
  assign new_n242_ = pi099 & pi104 & pi102 & pi103;
  assign new_n243_ = pi102 & pi107 & pi106 & pi105 & pi099;
  assign new_n244_ = new_n206_ | new_n236_ | new_n237_ | new_n235_;
  assign new_n245_ = new_n207_ | new_n239_ | new_n240_ | new_n238_;
  assign new_n246_ = new_n208_ | new_n242_ | new_n243_ | new_n241_;
  assign new_n247_ = pi110 & pi108 & pi109;
  assign new_n248_ = pi108 & pi113 & pi111 & pi112;
  assign new_n249_ = pi111 & pi116 & pi115 & pi114 & pi108;
  assign new_n250_ = pi119 & pi117 & pi118;
  assign new_n251_ = pi117 & pi122 & pi120 & pi121;
  assign new_n252_ = pi120 & pi125 & pi124 & pi123 & pi117;
  assign new_n253_ = pi128 & pi126 & pi127;
  assign new_n254_ = pi126 & pi131 & pi129 & pi130;
  assign new_n255_ = pi129 & pi134 & pi133 & pi132 & pi126;
  assign new_n256_ = pi137 & pi135 & pi136;
  assign new_n257_ = pi135 & pi140 & pi138 & pi139;
  assign new_n258_ = pi138 & pi143 & pi142 & pi141 & pi135;
  assign new_n259_ = new_n210_ | new_n251_ | new_n252_ | new_n250_;
  assign new_n260_ = new_n211_ | new_n254_ | new_n255_ | new_n253_;
  assign new_n261_ = new_n212_ | new_n257_ | new_n258_ | new_n256_;
  assign new_n262_ = pi146 & pi144 & pi145;
  assign new_n263_ = pi144 & pi149 & pi147 & pi148;
  assign new_n264_ = pi147 & pi152 & pi151 & pi150 & pi144;
  assign new_n265_ = pi155 & pi153 & pi154;
  assign new_n266_ = pi153 & pi158 & pi156 & pi157;
  assign new_n267_ = pi156 & pi161 & pi160 & pi159 & pi153;
  assign new_n268_ = pi164 & pi162 & pi163;
  assign new_n269_ = pi162 & pi167 & pi165 & pi166;
  assign new_n270_ = pi165 & pi170 & pi169 & pi168 & pi162;
  assign new_n271_ = pi173 & pi171 & pi172;
  assign new_n272_ = pi171 & pi176 & pi174 & pi175;
  assign new_n273_ = pi174 & pi179 & pi178 & pi177 & pi171;
  assign new_n274_ = new_n214_ | new_n266_ | new_n267_ | new_n265_;
  assign new_n275_ = new_n215_ | new_n269_ | new_n270_ | new_n268_;
  assign new_n276_ = new_n216_ | new_n272_ | new_n273_ | new_n271_;
  assign new_n277_ = pi180 & new_n229_;
  assign new_n278_ = pi180 & pi181 & new_n230_;
  assign new_n279_ = pi181 & new_n231_ & pi182 & pi180;
  assign new_n280_ = pi183 & new_n244_;
  assign new_n281_ = pi183 & pi184 & new_n245_;
  assign new_n282_ = pi184 & new_n246_ & pi185 & pi183;
  assign new_n283_ = pi186 & new_n259_;
  assign new_n284_ = pi186 & pi187 & new_n260_;
  assign new_n285_ = pi187 & new_n261_ & pi188 & pi186;
  assign new_n286_ = pi189 & new_n274_;
  assign new_n287_ = pi189 & pi190 & new_n275_;
  assign new_n288_ = pi190 & new_n276_ & pi191 & pi189;
  assign po2 = new_n218_ | new_n201_ | new_n279_ | new_n277_ | new_n278_ | new_n217_ | new_n219_;
  assign po3 = new_n233_ | new_n205_ | new_n282_ | new_n280_ | new_n281_ | new_n232_ | new_n234_;
  assign po4 = new_n248_ | new_n209_ | new_n285_ | new_n283_ | new_n284_ | new_n247_ | new_n249_;
  assign po5 = new_n263_ | new_n213_ | new_n288_ | new_n286_ | new_n287_ | new_n262_ | new_n264_;
endmodule


