// Benchmark "i2" written by ABC on Thu Mar 19 13:02:36 2020

module i2 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200,
    po0  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200;
  output po0;
  wire new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_;
  assign new_n203_ = pi030 | pi031 | pi028 | pi029 | pi026 | pi027 | pi024 | pi025 | pi022 | pi023 | pi020 | pi021 | pi018 | pi019 | pi016 | pi017 | pi014 | pi015 | pi012 | pi013 | pi010 | pi011 | pi008 | pi009 | pi006 | pi007 | pi004 | pi005 | pi002 | pi003 | pi000 | pi001;
  assign new_n204_ = pi062 | pi063 | pi060 | pi061 | pi058 | pi059 | pi056 | pi057 | pi054 | pi055 | pi052 | pi053 | pi050 | pi051 | pi048 | pi049 | pi046 | pi047 | pi044 | pi045 | pi042 | pi043 | pi040 | pi041 | pi038 | pi039 | pi036 | pi037 | pi034 | pi035 | pi032 | pi033;
  assign new_n205_ = pi094 | pi095 | pi092 | pi093 | pi090 | pi091 | pi088 | pi089 | pi086 | pi087 | pi084 | pi085 | pi082 | pi083 | pi080 | pi081 | pi078 | pi079 | pi076 | pi077 | pi074 | pi075 | pi072 | pi073 | pi070 | pi071 | pi068 | pi069 | pi066 | pi067 | pi064 | pi065;
  assign new_n206_ = pi126 | pi127 | pi124 | pi125 | pi122 | pi123 | pi120 | pi121 | pi118 | pi119 | pi116 | pi117 | pi114 | pi115 | pi112 | pi113 | pi110 | pi111 | pi108 | pi109 | pi106 | pi107 | pi104 | pi105 | pi102 | pi103 | pi100 | pi101 | pi098 | pi099 | pi096 | pi097;
  assign new_n207_ = ~pi128;
  assign new_n208_ = new_n207_ & pi129;
  assign new_n209_ = new_n207_ & pi130 & new_n203_;
  assign new_n210_ = new_n207_ & pi130 & new_n204_;
  assign new_n211_ = pi128 & pi131;
  assign new_n212_ = pi128 & pi130 & new_n205_;
  assign new_n213_ = pi128 & pi130 & new_n206_;
  assign new_n214_ = pi146 | pi147 | pi144 | pi145 | pi142 | pi143 | pi140 | pi141 | pi138 | pi139 | pi136 | pi137 | pi134 | pi135 | pi132 | pi133;
  assign new_n215_ = pi162 | pi163 | pi160 | pi161 | pi158 | pi159 | pi156 | pi157 | pi154 | pi155 | pi152 | pi153 | pi150 | pi151 | pi148 | pi149;
  assign new_n216_ = pi178 | pi179 | pi176 | pi177 | pi174 | pi175 | pi172 | pi173 | pi170 | pi171 | pi168 | pi169 | pi166 | pi167 | pi164 | pi165;
  assign new_n217_ = pi181 & pi180 & new_n214_;
  assign new_n218_ = pi181 & new_n215_;
  assign new_n219_ = pi180 & new_n218_;
  assign new_n220_ = pi181 & new_n216_;
  assign new_n221_ = pi180 & new_n220_;
  assign new_n222_ = pi180 & new_n216_;
  assign new_n223_ = pi184 | pi185 | pi182 | pi183;
  assign new_n224_ = pi188 | pi189 | pi186 | pi187;
  assign new_n225_ = pi192 | pi193 | pi190 | pi191;
  assign new_n226_ = pi195 & pi194 & new_n223_;
  assign new_n227_ = pi195 & new_n224_;
  assign new_n228_ = pi194 & new_n227_;
  assign new_n229_ = pi195 & new_n225_;
  assign new_n230_ = pi194 & new_n229_;
  assign new_n231_ = pi194 & new_n225_;
  assign new_n232_ = pi198 & pi196 & pi197;
  assign new_n233_ = pi198 & pi199;
  assign new_n234_ = pi196 & new_n233_;
  assign new_n235_ = pi198 & pi200;
  assign new_n236_ = pi196 & new_n235_;
  assign new_n237_ = pi196 & pi200;
  assign po0 = new_n235_ | new_n232_ | new_n236_ | new_n229_ | new_n226_ | new_n230_ | new_n220_ | new_n217_ | new_n221_ | new_n212_ | new_n208_ | new_n210_ | new_n209_ | new_n213_ | new_n211_ | new_n219_ | new_n222_ | new_n218_ | new_n228_ | new_n231_ | new_n227_ | new_n234_ | new_n237_ | new_n233_;
endmodule


