// Benchmark "t481" written by ABC on Thu Mar 19 13:02:36 2020

module t481 ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15,
    po0  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15;
  output po0;
  wire new_n18_, new_n19_, new_n20_, new_n21_, new_n22_, new_n23_, new_n24_,
    new_n25_, new_n26_, new_n27_, new_n28_, new_n29_, new_n30_, new_n31_,
    new_n32_, new_n33_, new_n34_, new_n35_, new_n36_, new_n37_, new_n38_,
    new_n39_, new_n40_, new_n41_, new_n42_, new_n43_, new_n44_, new_n45_,
    new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_, new_n52_,
    new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_, new_n59_,
    new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_, new_n66_,
    new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_, new_n73_,
    new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_,
    new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_,
    new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_,
    new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_, new_n111_, new_n112_, new_n113_,
    new_n114_, new_n115_, new_n116_, new_n117_, new_n118_, new_n119_,
    new_n120_, new_n121_, new_n122_, new_n123_, new_n124_, new_n125_,
    new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_,
    new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_,
    new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_,
    new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_,
    new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_,
    new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_,
    new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_,
    new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_,
    new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_,
    new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_,
    new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_,
    new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_,
    new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_,
    new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_,
    new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_,
    new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_,
    new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_,
    new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_,
    new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_,
    new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_,
    new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_,
    new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_,
    new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_,
    new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_,
    new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_,
    new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_,
    new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_,
    new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_,
    new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_,
    new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_,
    new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_,
    new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_,
    new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_,
    new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_,
    new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_,
    new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_,
    new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_,
    new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_,
    new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_,
    new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_,
    new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_,
    new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_,
    new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_,
    new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_,
    new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_,
    new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_,
    new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_,
    new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_,
    new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_,
    new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_,
    new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_,
    new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_,
    new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_,
    new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_,
    new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_,
    new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_,
    new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_,
    new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_,
    new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_,
    new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_,
    new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_,
    new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_,
    new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_,
    new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_,
    new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_,
    new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_,
    new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_,
    new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_,
    new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_,
    new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_,
    new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_,
    new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_,
    new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_,
    new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_,
    new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_,
    new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_,
    new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_,
    new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_,
    new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_,
    new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_,
    new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_,
    new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_,
    new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_,
    new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_,
    new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_,
    new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_,
    new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_,
    new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_,
    new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_,
    new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_,
    new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_,
    new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_,
    new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_,
    new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_,
    new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_,
    new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_,
    new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_,
    new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_,
    new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_,
    new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_,
    new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_,
    new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_,
    new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_,
    new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_,
    new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_,
    new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_,
    new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_,
    new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_,
    new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_,
    new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_,
    new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_,
    new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_,
    new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_,
    new_n1944_, new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_,
    new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_,
    new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_,
    new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_,
    new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_,
    new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_,
    new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_,
    new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_,
    new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_,
    new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_,
    new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_,
    new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_,
    new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_,
    new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_,
    new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_,
    new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_,
    new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_,
    new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_,
    new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_,
    new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_,
    new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_,
    new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_,
    new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_,
    new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_,
    new_n2088_;
  assign new_n18_ = ~pi02 & ~pi08 & ~pi01;
  assign new_n19_ = ~pi10;
  assign new_n20_ = ~pi09 | ~new_n18_ | ~new_n19_;
  assign new_n21_ = ~pi02 & ~pi09 & ~pi01;
  assign new_n22_ = ~pi11;
  assign new_n23_ = ~pi10 | ~new_n21_ | ~new_n22_;
  assign new_n24_ = ~pi01;
  assign new_n25_ = ~pi02;
  assign new_n26_ = ~pi13;
  assign new_n27_ = ~pi14;
  assign new_n28_ = ~new_n24_ | ~new_n25_ | ~new_n26_ | ~new_n27_;
  assign new_n29_ = ~new_n24_ | ~new_n25_ | ~new_n26_ | ~pi15;
  assign new_n30_ = ~new_n20_ | ~new_n23_ | ~new_n28_ | ~new_n29_;
  assign new_n31_ = ~pi01 & ~pi02;
  assign new_n32_ = ~pi08 | ~new_n31_ | ~new_n22_ | ~pi10;
  assign new_n33_ = ~pi02 & ~pi08 & ~pi01;
  assign new_n34_ = ~pi11 | ~new_n33_ | ~pi09;
  assign new_n35_ = ~new_n24_ | ~new_n25_ | ~pi15 | ~pi12;
  assign new_n36_ = ~pi02 & ~pi12 & ~pi01;
  assign new_n37_ = ~pi15;
  assign new_n38_ = ~new_n36_ | ~new_n37_ | ~pi13 | ~pi14;
  assign new_n39_ = ~new_n32_ | ~new_n34_ | ~new_n35_ | ~new_n38_;
  assign new_n40_ = ~new_n24_ | ~new_n25_ | ~new_n27_ | ~pi12;
  assign new_n41_ = ~pi00;
  assign new_n42_ = ~new_n41_ & ~pi08 & ~pi02;
  assign new_n43_ = ~pi09 | ~new_n42_ | ~new_n19_;
  assign new_n44_ = ~new_n41_ & ~pi09 & ~pi02;
  assign new_n45_ = ~pi10 | ~new_n44_ | ~new_n22_;
  assign new_n46_ = ~new_n25_ | ~pi00 | ~new_n26_ | ~new_n27_;
  assign new_n47_ = ~new_n40_ | ~new_n43_ | ~new_n45_ | ~new_n46_;
  assign new_n48_ = ~new_n25_ | ~pi00 | ~new_n26_ | ~pi15;
  assign new_n49_ = ~pi11 & ~new_n19_;
  assign new_n50_ = ~new_n49_ | ~pi08 | ~new_n25_ | ~pi00;
  assign new_n51_ = ~new_n41_ & ~pi08 & ~pi02;
  assign new_n52_ = ~pi11 | ~new_n51_ | ~pi09;
  assign new_n53_ = ~new_n25_ | ~pi00 | ~pi15 | ~pi12;
  assign new_n54_ = ~new_n48_ | ~new_n50_ | ~new_n52_ | ~new_n53_;
  assign new_n55_ = ~new_n54_ & ~new_n47_ & ~new_n30_ & ~new_n39_;
  assign new_n56_ = ~pi04;
  assign new_n57_ = ~pi06;
  assign new_n58_ = ~new_n57_ & ~pi07 & ~new_n56_;
  assign new_n59_ = ~pi12 | ~new_n58_ | ~pi15;
  assign new_n60_ = ~pi12 & ~pi07 & ~new_n56_ & ~new_n57_;
  assign new_n61_ = ~new_n60_ | ~new_n37_ | ~pi13 | ~pi14;
  assign new_n62_ = ~pi12;
  assign new_n63_ = ~pi14 & ~new_n62_;
  assign new_n64_ = ~pi07;
  assign new_n65_ = ~new_n63_ | ~new_n64_ | ~pi04 | ~pi06;
  assign new_n66_ = ~pi03;
  assign new_n67_ = ~new_n66_ & ~pi08 & ~pi01;
  assign new_n68_ = ~pi09 | ~new_n67_ | ~new_n19_;
  assign new_n69_ = ~new_n59_ | ~new_n61_ | ~new_n65_ | ~new_n68_;
  assign new_n70_ = ~new_n37_ & ~pi13 & ~pi01 & ~new_n66_;
  assign new_n71_ = ~new_n22_ | ~pi10;
  assign new_n72_ = ~new_n66_ & ~pi01 & ~new_n71_ & ~pi09;
  assign new_n73_ = ~pi14 & ~pi13 & ~pi01 & ~new_n66_;
  assign new_n74_ = ~new_n73_ & ~new_n72_ & ~new_n69_ & ~new_n70_;
  assign new_n75_ = ~pi14 | ~new_n37_ | ~pi13;
  assign new_n76_ = ~new_n41_ & ~pi02 & ~new_n75_ & ~pi12;
  assign new_n77_ = ~new_n62_ & ~pi14 & ~pi02 & ~new_n41_;
  assign new_n78_ = ~pi06 | ~new_n64_ | ~pi04;
  assign new_n79_ = ~pi09;
  assign new_n80_ = ~new_n79_ & ~pi08 & ~new_n78_ & ~pi10;
  assign new_n81_ = ~pi06 | ~new_n64_ | ~pi04;
  assign new_n82_ = ~new_n19_ & ~pi09 & ~new_n81_ & ~pi11;
  assign new_n83_ = ~new_n82_ & ~new_n80_ & ~new_n76_ & ~new_n77_;
  assign new_n84_ = ~pi04 | ~pi06;
  assign new_n85_ = ~pi14 & ~pi13 & ~pi07 & ~new_n84_;
  assign new_n86_ = ~pi04 | ~pi06;
  assign new_n87_ = ~new_n37_ & ~pi13 & ~pi07 & ~new_n86_;
  assign new_n88_ = ~pi06 | ~new_n64_ | ~pi04;
  assign new_n89_ = ~pi08;
  assign new_n90_ = ~new_n19_ & ~new_n89_ & ~new_n88_ & ~pi11;
  assign new_n91_ = ~pi06 | ~new_n64_ | ~pi04;
  assign new_n92_ = ~new_n79_ & ~pi08 & ~new_n91_ & ~new_n22_;
  assign new_n93_ = ~new_n92_ & ~new_n90_ & ~new_n85_ & ~new_n87_;
  assign new_n94_ = ~new_n55_ | ~new_n74_ | ~new_n83_ | ~new_n93_;
  assign new_n95_ = ~pi05 | ~new_n57_ | ~new_n56_;
  assign new_n96_ = ~new_n79_ & ~pi08 & ~new_n95_ & ~pi10;
  assign new_n97_ = ~pi05 | ~new_n57_ | ~new_n56_;
  assign new_n98_ = ~new_n19_ & ~pi09 & ~new_n97_ & ~pi11;
  assign new_n99_ = ~new_n56_ | ~pi05;
  assign new_n100_ = ~pi14 & ~pi13 & ~pi06 & ~new_n99_;
  assign new_n101_ = ~new_n56_ | ~pi05;
  assign new_n102_ = ~new_n37_ & ~pi13 & ~pi06 & ~new_n101_;
  assign new_n103_ = ~new_n102_ & ~new_n100_ & ~new_n96_ & ~new_n98_;
  assign new_n104_ = ~pi05;
  assign new_n105_ = ~new_n104_ & ~pi06 & ~pi04;
  assign new_n106_ = ~pi12 | ~new_n105_ | ~pi15;
  assign new_n107_ = ~new_n104_ & ~pi06 & ~pi04;
  assign new_n108_ = ~new_n107_ | ~new_n22_ | ~pi08 | ~pi10;
  assign new_n109_ = ~new_n104_ & ~pi06 & ~pi04;
  assign new_n110_ = ~new_n109_ | ~pi11 | ~new_n89_ | ~pi09;
  assign new_n111_ = ~new_n103_ | ~new_n106_ | ~new_n108_ | ~new_n110_;
  assign new_n112_ = ~new_n57_ & ~pi07 & ~pi05;
  assign new_n113_ = ~new_n112_ | ~new_n22_ | ~new_n79_ | ~pi10;
  assign new_n114_ = ~pi13 & ~pi14;
  assign new_n115_ = ~new_n114_ | ~new_n64_ | ~new_n104_ | ~pi06;
  assign new_n116_ = ~new_n57_ & ~pi07 & ~pi05;
  assign new_n117_ = ~pi15 | ~new_n116_ | ~new_n26_;
  assign new_n118_ = ~new_n57_ & ~pi07 & ~pi05;
  assign new_n119_ = ~new_n118_ | ~new_n22_ | ~pi08 | ~pi10;
  assign new_n120_ = ~new_n113_ | ~new_n115_ | ~new_n117_ | ~new_n119_;
  assign new_n121_ = ~new_n57_ & ~pi07 & ~pi05;
  assign new_n122_ = ~new_n121_ | ~pi11 | ~new_n89_ | ~pi09;
  assign new_n123_ = ~new_n57_ & ~pi07 & ~pi05;
  assign new_n124_ = ~pi12 | ~new_n123_ | ~pi15;
  assign new_n125_ = ~pi12 & ~pi07 & ~pi05 & ~new_n57_;
  assign new_n126_ = ~new_n125_ | ~new_n37_ | ~pi13 | ~pi14;
  assign new_n127_ = ~new_n57_ & ~pi07 & ~pi05;
  assign new_n128_ = ~pi12 | ~new_n127_ | ~new_n27_;
  assign new_n129_ = ~new_n122_ | ~new_n124_ | ~new_n126_ | ~new_n128_;
  assign new_n130_ = ~new_n129_ & ~new_n111_ & ~new_n120_;
  assign new_n131_ = ~pi00 | ~pi03 | ~new_n26_ | ~pi15;
  assign new_n132_ = ~pi11 & ~new_n19_;
  assign new_n133_ = ~new_n132_ | ~pi08 | ~pi00 | ~pi03;
  assign new_n134_ = ~new_n66_ & ~pi08 & ~new_n41_;
  assign new_n135_ = ~pi11 | ~new_n134_ | ~pi09;
  assign new_n136_ = ~pi00 | ~pi03 | ~pi15 | ~pi12;
  assign new_n137_ = ~new_n131_ | ~new_n133_ | ~new_n135_ | ~new_n136_;
  assign new_n138_ = ~pi06 | ~new_n64_ | ~new_n104_;
  assign new_n139_ = ~new_n79_ & ~pi08 & ~new_n138_ & ~pi10;
  assign new_n140_ = ~pi03 | ~new_n62_ | ~pi00;
  assign new_n141_ = ~new_n27_ & ~new_n26_ & ~new_n140_ & ~pi15;
  assign new_n142_ = ~new_n62_ & ~pi14 & ~new_n41_ & ~new_n66_;
  assign new_n143_ = ~new_n142_ & ~new_n141_ & ~new_n137_ & ~new_n139_;
  assign new_n144_ = ~pi03 | ~pi08 | ~new_n24_;
  assign new_n145_ = ~new_n19_ & ~new_n144_ & ~pi11;
  assign new_n146_ = ~pi09 | ~pi11;
  assign new_n147_ = ~new_n66_ & ~pi01 & ~new_n146_ & ~pi08;
  assign new_n148_ = ~new_n62_ & ~new_n37_ & ~pi01 & ~new_n66_;
  assign new_n149_ = ~pi14 | ~new_n37_ | ~pi13;
  assign new_n150_ = ~new_n66_ & ~pi01 & ~new_n149_ & ~pi12;
  assign new_n151_ = ~new_n150_ & ~new_n148_ & ~new_n145_ & ~new_n147_;
  assign new_n152_ = ~new_n62_ & ~pi14 & ~pi01 & ~new_n66_;
  assign new_n153_ = ~pi00 | ~pi03;
  assign new_n154_ = ~new_n79_ & ~pi10 & ~pi08 & ~new_n153_;
  assign new_n155_ = ~pi00 | ~pi03;
  assign new_n156_ = ~new_n19_ & ~pi11 & ~pi09 & ~new_n155_;
  assign new_n157_ = ~pi14 & ~pi13 & ~new_n41_ & ~new_n66_;
  assign new_n158_ = ~new_n157_ & ~new_n156_ & ~new_n152_ & ~new_n154_;
  assign new_n159_ = ~new_n130_ | ~new_n143_ | ~new_n151_ | ~new_n158_;
  assign new_n160_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n161_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n162_ = ~pi08 | ~pi11 | ~new_n64_;
  assign new_n163_ = ~pi12 | ~new_n37_ | ~pi14;
  assign new_n164_ = ~new_n163_ & ~new_n162_ & ~new_n160_ & ~new_n161_;
  assign new_n165_ = ~pi05 & ~pi06;
  assign new_n166_ = ~new_n165_ | ~new_n25_ | ~new_n41_ | ~pi01;
  assign new_n167_ = ~pi11 | ~pi12 | ~pi08;
  assign new_n168_ = ~new_n27_ & ~pi15 & ~new_n166_ & ~new_n167_;
  assign new_n169_ = ~pi05 & ~pi06;
  assign new_n170_ = ~new_n169_ | ~pi03 | ~new_n41_ | ~pi01;
  assign new_n171_ = ~pi11 | ~pi12 | ~pi08;
  assign new_n172_ = ~new_n27_ & ~pi15 & ~new_n170_ & ~new_n171_;
  assign new_n173_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n174_ = ~pi04 | ~new_n173_ | ~new_n57_;
  assign new_n175_ = ~pi11 | ~pi12 | ~pi08;
  assign new_n176_ = ~new_n27_ & ~pi15 & ~new_n174_ & ~new_n175_;
  assign new_n177_ = ~new_n176_ & ~new_n172_ & ~new_n164_ & ~new_n168_;
  assign new_n178_ = ~pi11 | ~pi12 | ~pi08;
  assign new_n179_ = ~new_n27_ & ~new_n178_ & ~pi15;
  assign new_n180_ = ~new_n24_ & ~new_n66_ & ~pi00;
  assign new_n181_ = ~new_n179_ | ~new_n180_ | ~new_n104_ | ~pi07;
  assign new_n182_ = ~pi11 | ~pi12 | ~pi08;
  assign new_n183_ = ~new_n27_ & ~new_n182_ & ~pi15;
  assign new_n184_ = ~new_n24_ & ~new_n66_ & ~pi00;
  assign new_n185_ = ~new_n183_ | ~new_n184_ | ~new_n57_ | ~pi04;
  assign new_n186_ = ~pi11 | ~pi12 | ~pi08;
  assign new_n187_ = ~new_n27_ & ~new_n186_ & ~pi15;
  assign new_n188_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n189_ = ~new_n187_ | ~new_n188_ | ~new_n104_ | ~pi07;
  assign new_n190_ = ~new_n177_ | ~new_n181_ | ~new_n185_ | ~new_n189_;
  assign new_n191_ = ~new_n25_ & ~pi03 & ~pi00 & ~new_n24_;
  assign new_n192_ = ~new_n191_ | ~new_n22_ | ~pi08 | ~pi10;
  assign new_n193_ = ~new_n25_ & ~pi03 & ~pi00 & ~new_n24_;
  assign new_n194_ = ~new_n193_ | ~pi11 | ~new_n89_ | ~pi09;
  assign new_n195_ = ~new_n24_ & ~new_n25_ & ~pi00;
  assign new_n196_ = ~new_n195_ | ~pi15 | ~new_n66_ | ~pi12;
  assign new_n197_ = ~new_n25_ & ~pi03 & ~pi00 & ~new_n24_;
  assign new_n198_ = ~new_n27_ & ~pi15 & ~pi12 & ~new_n26_;
  assign new_n199_ = ~new_n197_ | ~new_n198_;
  assign new_n200_ = ~new_n192_ | ~new_n194_ | ~new_n196_ | ~new_n199_;
  assign new_n201_ = ~new_n62_ & ~pi14 & ~pi03;
  assign new_n202_ = ~new_n201_ | ~pi02 | ~new_n41_ | ~pi01;
  assign new_n203_ = ~pi11 | ~pi12 | ~pi08;
  assign new_n204_ = ~new_n27_ & ~new_n203_ & ~pi15;
  assign new_n205_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n206_ = ~new_n204_ | ~new_n205_ | ~pi07 | ~pi04;
  assign new_n207_ = ~pi11 | ~pi12 | ~pi08;
  assign new_n208_ = ~new_n27_ & ~new_n207_ & ~pi15;
  assign new_n209_ = ~new_n24_ & ~new_n66_ & ~pi00;
  assign new_n210_ = ~new_n208_ | ~new_n209_ | ~pi07 | ~pi04;
  assign new_n211_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n212_ = ~new_n24_ & ~pi00 & ~new_n211_ & ~pi02;
  assign new_n213_ = ~pi08 | ~pi11 | ~new_n64_;
  assign new_n214_ = ~new_n62_ & ~new_n27_ & ~new_n213_ & ~pi15;
  assign new_n215_ = ~new_n212_ | ~new_n214_;
  assign new_n216_ = ~new_n202_ | ~new_n206_ | ~new_n210_ | ~new_n215_;
  assign new_n217_ = ~new_n216_ & ~new_n190_ & ~new_n200_;
  assign new_n218_ = ~pi04 & ~new_n104_;
  assign new_n219_ = ~pi07 | ~new_n218_ | ~pi15 | ~pi12;
  assign new_n220_ = ~new_n64_ & ~pi12 & ~pi04 & ~new_n104_;
  assign new_n221_ = ~new_n220_ | ~new_n37_ | ~pi13 | ~pi14;
  assign new_n222_ = ~pi04 & ~new_n104_;
  assign new_n223_ = ~pi07 | ~new_n222_ | ~new_n27_ | ~pi12;
  assign new_n224_ = ~new_n25_ & ~pi03 & ~pi00 & ~new_n24_;
  assign new_n225_ = ~new_n224_ | ~new_n19_ | ~new_n89_ | ~pi09;
  assign new_n226_ = ~new_n219_ | ~new_n221_ | ~new_n223_ | ~new_n225_;
  assign new_n227_ = ~pi01 | ~pi02 | ~new_n41_;
  assign new_n228_ = ~pi13 & ~pi03 & ~new_n227_ & ~new_n37_;
  assign new_n229_ = ~new_n41_ | ~pi01 | ~new_n66_ | ~pi02;
  assign new_n230_ = ~new_n19_ & ~pi09 & ~new_n229_ & ~pi11;
  assign new_n231_ = ~pi01 | ~pi02 | ~new_n41_;
  assign new_n232_ = ~pi13 & ~pi03 & ~new_n231_ & ~pi14;
  assign new_n233_ = ~new_n232_ & ~new_n230_ & ~new_n226_ & ~new_n228_;
  assign new_n234_ = ~new_n56_ | ~pi05 | ~new_n57_ | ~new_n62_;
  assign new_n235_ = ~new_n27_ & ~new_n26_ & ~new_n234_ & ~pi15;
  assign new_n236_ = ~new_n56_ | ~pi05;
  assign new_n237_ = ~new_n62_ & ~pi14 & ~pi06 & ~new_n236_;
  assign new_n238_ = ~pi05 | ~pi07 | ~new_n56_;
  assign new_n239_ = ~new_n79_ & ~pi08 & ~new_n238_ & ~pi10;
  assign new_n240_ = ~pi05 | ~pi07 | ~new_n56_;
  assign new_n241_ = ~new_n19_ & ~pi09 & ~new_n240_ & ~pi11;
  assign new_n242_ = ~new_n241_ & ~new_n239_ & ~new_n235_ & ~new_n237_;
  assign new_n243_ = ~pi05 | ~pi07 | ~new_n56_;
  assign new_n244_ = ~pi14 & ~new_n243_ & ~pi13;
  assign new_n245_ = ~pi05 | ~pi07 | ~new_n56_;
  assign new_n246_ = ~new_n37_ & ~new_n245_ & ~pi13;
  assign new_n247_ = ~pi05 | ~pi07 | ~new_n56_;
  assign new_n248_ = ~new_n19_ & ~new_n89_ & ~new_n247_ & ~pi11;
  assign new_n249_ = ~pi05 | ~pi07 | ~new_n56_;
  assign new_n250_ = ~new_n79_ & ~pi08 & ~new_n249_ & ~new_n22_;
  assign new_n251_ = ~new_n250_ & ~new_n248_ & ~new_n244_ & ~new_n246_;
  assign new_n252_ = ~new_n217_ | ~new_n233_ | ~new_n242_ | ~new_n251_;
  assign new_n253_ = ~pi06 & ~new_n56_;
  assign new_n254_ = ~new_n253_ | ~new_n66_ | ~pi02 | ~pi00;
  assign new_n255_ = ~pi08 | ~pi12 | ~new_n19_;
  assign new_n256_ = ~new_n27_ & ~pi15 & ~new_n254_ & ~new_n255_;
  assign new_n257_ = ~new_n89_ & ~pi10 & ~pi07;
  assign new_n258_ = ~new_n257_ | ~new_n37_ | ~pi14 | ~pi12;
  assign new_n259_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n260_ = ~new_n24_ | ~pi02;
  assign new_n261_ = ~new_n260_ & ~pi03 & ~new_n258_ & ~new_n259_;
  assign new_n262_ = ~new_n89_ & ~pi10 & ~pi07;
  assign new_n263_ = ~new_n262_ | ~new_n37_ | ~pi14 | ~pi12;
  assign new_n264_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n265_ = ~pi02 | ~pi00;
  assign new_n266_ = ~new_n265_ & ~pi03 & ~new_n263_ & ~new_n264_;
  assign new_n267_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n268_ = ~pi07 | ~new_n267_ | ~new_n104_;
  assign new_n269_ = ~pi08 | ~pi12 | ~new_n19_;
  assign new_n270_ = ~new_n27_ & ~pi15 & ~new_n268_ & ~new_n269_;
  assign new_n271_ = ~new_n270_ & ~new_n266_ & ~new_n256_ & ~new_n261_;
  assign new_n272_ = ~pi08 | ~pi12 | ~new_n19_;
  assign new_n273_ = ~new_n27_ & ~new_n272_ & ~pi15;
  assign new_n274_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n275_ = ~new_n273_ | ~new_n274_ | ~pi07 | ~pi04;
  assign new_n276_ = ~pi02 | ~pi00;
  assign new_n277_ = ~new_n64_ & ~pi05 & ~pi03 & ~new_n276_;
  assign new_n278_ = ~new_n89_ & ~new_n62_ & ~pi10;
  assign new_n279_ = ~new_n277_ | ~new_n278_ | ~new_n37_ | ~pi14;
  assign new_n280_ = ~pi07 | ~pi04;
  assign new_n281_ = ~new_n24_ & ~pi00 & ~new_n280_ & ~pi02;
  assign new_n282_ = ~pi10 & ~new_n62_ & ~pi09;
  assign new_n283_ = ~new_n281_ | ~new_n282_ | ~new_n37_ | ~pi14;
  assign new_n284_ = ~new_n271_ | ~new_n275_ | ~new_n279_ | ~new_n283_;
  assign new_n285_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n286_ = ~pi06 & ~new_n285_ & ~pi05;
  assign new_n287_ = ~new_n89_ & ~new_n62_ & ~pi10;
  assign new_n288_ = ~new_n286_ | ~new_n287_ | ~new_n37_ | ~pi14;
  assign new_n289_ = ~pi08 | ~pi12 | ~new_n19_;
  assign new_n290_ = ~new_n27_ & ~new_n289_ & ~pi15;
  assign new_n291_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n292_ = ~new_n290_ | ~new_n291_ | ~new_n57_ | ~pi04;
  assign new_n293_ = ~pi08 | ~pi12 | ~new_n19_;
  assign new_n294_ = ~new_n27_ & ~new_n293_ & ~pi15;
  assign new_n295_ = ~new_n24_ & ~new_n66_ & ~pi00;
  assign new_n296_ = ~new_n294_ | ~new_n295_ | ~new_n57_ | ~pi04;
  assign new_n297_ = ~pi08 | ~pi12 | ~new_n19_;
  assign new_n298_ = ~new_n27_ & ~new_n297_ & ~pi15;
  assign new_n299_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n300_ = ~new_n298_ | ~new_n299_ | ~new_n104_ | ~pi07;
  assign new_n301_ = ~new_n288_ | ~new_n292_ | ~new_n296_ | ~new_n300_;
  assign new_n302_ = ~pi08 | ~pi12 | ~new_n19_;
  assign new_n303_ = ~new_n27_ & ~new_n302_ & ~pi15;
  assign new_n304_ = ~new_n24_ & ~new_n66_ & ~pi00;
  assign new_n305_ = ~new_n303_ | ~new_n304_ | ~new_n104_ | ~pi07;
  assign new_n306_ = ~new_n24_ | ~pi02;
  assign new_n307_ = ~pi06 & ~pi05 & ~pi03 & ~new_n306_;
  assign new_n308_ = ~new_n89_ & ~new_n62_ & ~pi10;
  assign new_n309_ = ~new_n307_ | ~new_n308_ | ~new_n37_ | ~pi14;
  assign new_n310_ = ~pi02 | ~pi00;
  assign new_n311_ = ~pi06 & ~pi05 & ~pi03 & ~new_n310_;
  assign new_n312_ = ~new_n89_ & ~new_n62_ & ~pi10;
  assign new_n313_ = ~new_n311_ | ~new_n312_ | ~new_n37_ | ~pi14;
  assign new_n314_ = ~pi08 | ~pi12 | ~new_n19_;
  assign new_n315_ = ~new_n27_ & ~new_n314_ & ~pi15;
  assign new_n316_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n317_ = ~new_n315_ | ~new_n316_ | ~new_n57_ | ~pi04;
  assign new_n318_ = ~new_n305_ | ~new_n309_ | ~new_n313_ | ~new_n317_;
  assign new_n319_ = ~new_n318_ & ~new_n284_ & ~new_n301_;
  assign new_n320_ = ~pi08 | ~pi12 | ~new_n19_;
  assign new_n321_ = ~new_n27_ & ~new_n320_ & ~pi15;
  assign new_n322_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n323_ = ~new_n321_ | ~new_n322_ | ~pi07 | ~pi04;
  assign new_n324_ = ~pi11 | ~pi12 | ~pi08;
  assign new_n325_ = ~new_n27_ & ~new_n324_ & ~pi15;
  assign new_n326_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n327_ = ~new_n325_ | ~new_n326_ | ~pi07 | ~pi04;
  assign new_n328_ = ~pi11 | ~pi12 | ~pi08;
  assign new_n329_ = ~new_n27_ & ~new_n328_ & ~pi15;
  assign new_n330_ = ~new_n41_ & ~pi03 & ~new_n25_;
  assign new_n331_ = ~new_n329_ | ~new_n330_ | ~pi07 | ~pi04;
  assign new_n332_ = ~pi08 | ~pi12 | ~new_n19_;
  assign new_n333_ = ~new_n27_ & ~new_n332_ & ~pi15;
  assign new_n334_ = ~new_n24_ & ~new_n66_ & ~pi00;
  assign new_n335_ = ~new_n333_ | ~new_n334_ | ~pi07 | ~pi04;
  assign new_n336_ = ~new_n323_ | ~new_n327_ | ~new_n331_ | ~new_n335_;
  assign new_n337_ = ~pi05 & ~pi06;
  assign new_n338_ = ~new_n337_ | ~new_n25_ | ~new_n41_ | ~pi01;
  assign new_n339_ = ~pi08 | ~pi12 | ~new_n19_;
  assign new_n340_ = ~new_n27_ & ~pi15 & ~new_n338_ & ~new_n339_;
  assign new_n341_ = ~new_n89_ & ~pi10 & ~pi07;
  assign new_n342_ = ~new_n341_ | ~new_n37_ | ~pi14 | ~pi12;
  assign new_n343_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n344_ = ~new_n41_ | ~pi01;
  assign new_n345_ = ~new_n344_ & ~pi02 & ~new_n342_ & ~new_n343_;
  assign new_n346_ = ~new_n89_ & ~pi10 & ~pi07;
  assign new_n347_ = ~new_n346_ | ~new_n37_ | ~pi14 | ~pi12;
  assign new_n348_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n349_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n350_ = ~new_n349_ & ~new_n347_ & ~new_n348_;
  assign new_n351_ = ~new_n350_ & ~new_n345_ & ~new_n336_ & ~new_n340_;
  assign new_n352_ = ~pi05 & ~pi06;
  assign new_n353_ = ~new_n352_ | ~new_n66_ | ~new_n24_ | ~pi02;
  assign new_n354_ = ~pi11 | ~pi12 | ~pi08;
  assign new_n355_ = ~new_n27_ & ~pi15 & ~new_n353_ & ~new_n354_;
  assign new_n356_ = ~pi05 & ~pi06;
  assign new_n357_ = ~new_n356_ | ~new_n66_ | ~pi02 | ~pi00;
  assign new_n358_ = ~pi11 | ~pi12 | ~pi08;
  assign new_n359_ = ~new_n27_ & ~pi15 & ~new_n357_ & ~new_n358_;
  assign new_n360_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n361_ = ~pi04 | ~new_n360_ | ~new_n57_;
  assign new_n362_ = ~pi11 | ~pi12 | ~pi08;
  assign new_n363_ = ~new_n27_ & ~pi15 & ~new_n361_ & ~new_n362_;
  assign new_n364_ = ~pi06 & ~new_n56_;
  assign new_n365_ = ~new_n364_ | ~new_n66_ | ~pi02 | ~pi00;
  assign new_n366_ = ~pi11 | ~pi12 | ~pi08;
  assign new_n367_ = ~new_n27_ & ~pi15 & ~new_n365_ & ~new_n366_;
  assign new_n368_ = ~new_n367_ & ~new_n363_ & ~new_n355_ & ~new_n359_;
  assign new_n369_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n370_ = ~new_n369_ | ~pi06 | ~new_n56_ | ~pi05;
  assign new_n371_ = ~pi08 | ~pi11 | ~new_n64_;
  assign new_n372_ = ~pi14 | ~pi12;
  assign new_n373_ = ~new_n372_ & ~pi15 & ~new_n370_ & ~new_n371_;
  assign new_n374_ = ~pi00 | ~new_n66_ | ~pi02;
  assign new_n375_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n376_ = ~pi08 | ~pi11 | ~new_n64_;
  assign new_n377_ = ~pi12 | ~new_n37_ | ~pi14;
  assign new_n378_ = ~new_n377_ & ~new_n376_ & ~new_n374_ & ~new_n375_;
  assign new_n379_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n380_ = ~pi07 | ~new_n379_ | ~new_n104_;
  assign new_n381_ = ~pi11 | ~pi12 | ~pi08;
  assign new_n382_ = ~new_n27_ & ~pi15 & ~new_n380_ & ~new_n381_;
  assign new_n383_ = ~pi05 & ~new_n64_;
  assign new_n384_ = ~new_n383_ | ~new_n66_ | ~pi02 | ~pi00;
  assign new_n385_ = ~pi11 | ~pi12 | ~pi08;
  assign new_n386_ = ~new_n27_ & ~pi15 & ~new_n384_ & ~new_n385_;
  assign new_n387_ = ~new_n386_ & ~new_n382_ & ~new_n373_ & ~new_n378_;
  assign new_n388_ = ~new_n319_ | ~new_n351_ | ~new_n368_ | ~new_n387_;
  assign new_n389_ = ~new_n388_ & ~new_n252_ & ~new_n94_ & ~new_n159_;
  assign new_n390_ = ~pi12 | ~new_n37_ | ~pi14;
  assign new_n391_ = ~pi09 & ~pi07 & ~new_n390_ & ~pi10;
  assign new_n392_ = ~new_n41_ & ~pi03 & ~new_n25_;
  assign new_n393_ = ~pi04 & ~new_n104_;
  assign new_n394_ = ~new_n391_ | ~new_n392_ | ~pi06 | ~new_n393_;
  assign new_n395_ = ~new_n104_ | ~pi07;
  assign new_n396_ = ~new_n25_ & ~pi01 & ~new_n395_ & ~pi03;
  assign new_n397_ = ~pi10 & ~new_n62_ & ~pi09;
  assign new_n398_ = ~new_n396_ | ~new_n397_ | ~new_n37_ | ~pi14;
  assign new_n399_ = ~pi02 | ~pi00;
  assign new_n400_ = ~new_n64_ & ~pi05 & ~pi03 & ~new_n399_;
  assign new_n401_ = ~pi10 & ~new_n62_ & ~pi09;
  assign new_n402_ = ~new_n400_ | ~new_n401_ | ~new_n37_ | ~pi14;
  assign new_n403_ = ~pi07 | ~pi04;
  assign new_n404_ = ~new_n24_ & ~pi00 & ~new_n403_ & ~pi02;
  assign new_n405_ = ~pi10 & ~pi13 & ~pi09;
  assign new_n406_ = ~new_n404_ | ~new_n405_ | ~new_n37_ | ~pi14;
  assign new_n407_ = ~new_n394_ | ~new_n398_ | ~new_n402_ | ~new_n406_;
  assign new_n408_ = ~pi07 | ~pi04;
  assign new_n409_ = ~new_n25_ & ~pi01 & ~new_n408_ & ~pi03;
  assign new_n410_ = ~pi10 & ~new_n62_ & ~pi09;
  assign new_n411_ = ~new_n409_ | ~new_n410_ | ~new_n37_ | ~pi14;
  assign new_n412_ = ~pi07 | ~pi04;
  assign new_n413_ = ~new_n41_ & ~new_n25_ & ~new_n412_ & ~pi03;
  assign new_n414_ = ~pi10 & ~new_n62_ & ~pi09;
  assign new_n415_ = ~new_n413_ | ~new_n414_ | ~new_n37_ | ~pi14;
  assign new_n416_ = ~pi07 | ~pi04;
  assign new_n417_ = ~new_n24_ & ~pi00 & ~new_n416_ & ~new_n66_;
  assign new_n418_ = ~pi10 & ~pi13 & ~pi09;
  assign new_n419_ = ~new_n417_ | ~new_n418_ | ~new_n37_ | ~pi14;
  assign new_n420_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n421_ = ~new_n24_ & ~pi00 & ~new_n420_ & ~pi02;
  assign new_n422_ = ~pi09 & ~pi10 & ~pi07;
  assign new_n423_ = ~new_n27_ & ~pi15 & ~pi13;
  assign new_n424_ = ~new_n423_ | ~new_n421_ | ~new_n422_;
  assign new_n425_ = ~new_n411_ | ~new_n415_ | ~new_n419_ | ~new_n424_;
  assign new_n426_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n427_ = ~new_n24_ & ~pi00 & ~new_n426_ & ~new_n66_;
  assign new_n428_ = ~pi09 & ~pi10 & ~pi07;
  assign new_n429_ = ~new_n27_ & ~pi15 & ~pi13;
  assign new_n430_ = ~new_n429_ | ~new_n427_ | ~new_n428_;
  assign new_n431_ = ~new_n41_ | ~pi01;
  assign new_n432_ = ~pi06 & ~pi05 & ~pi02 & ~new_n431_;
  assign new_n433_ = ~pi10 & ~pi13 & ~pi09;
  assign new_n434_ = ~new_n432_ | ~new_n433_ | ~new_n37_ | ~pi14;
  assign new_n435_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n436_ = ~pi06 & ~new_n435_ & ~pi05;
  assign new_n437_ = ~pi10 & ~pi13 & ~pi09;
  assign new_n438_ = ~new_n436_ | ~new_n437_ | ~new_n37_ | ~pi14;
  assign new_n439_ = ~new_n57_ | ~pi04;
  assign new_n440_ = ~new_n24_ & ~pi00 & ~new_n439_ & ~pi02;
  assign new_n441_ = ~pi10 & ~pi13 & ~pi09;
  assign new_n442_ = ~new_n440_ | ~new_n441_ | ~new_n37_ | ~pi14;
  assign new_n443_ = ~new_n430_ | ~new_n434_ | ~new_n438_ | ~new_n442_;
  assign new_n444_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n445_ = ~new_n64_ & ~new_n444_ & ~pi05;
  assign new_n446_ = ~pi10 & ~pi13 & ~pi09;
  assign new_n447_ = ~new_n445_ | ~new_n446_ | ~new_n37_ | ~pi14;
  assign new_n448_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n449_ = ~new_n56_ & ~new_n448_ & ~pi06;
  assign new_n450_ = ~pi10 & ~pi13 & ~pi09;
  assign new_n451_ = ~new_n449_ | ~new_n450_ | ~new_n37_ | ~pi14;
  assign new_n452_ = ~new_n104_ | ~pi07;
  assign new_n453_ = ~new_n24_ & ~pi00 & ~new_n452_ & ~pi02;
  assign new_n454_ = ~pi10 & ~pi13 & ~pi09;
  assign new_n455_ = ~new_n453_ | ~new_n454_ | ~new_n37_ | ~pi14;
  assign new_n456_ = ~new_n455_ | ~new_n447_ | ~new_n451_;
  assign new_n457_ = ~new_n456_ & ~new_n443_ & ~new_n407_ & ~new_n425_;
  assign new_n458_ = ~new_n104_ | ~pi07;
  assign new_n459_ = ~new_n24_ & ~pi00 & ~new_n458_ & ~pi02;
  assign new_n460_ = ~pi10 & ~new_n62_ & ~pi09;
  assign new_n461_ = ~new_n459_ | ~new_n460_ | ~new_n37_ | ~pi14;
  assign new_n462_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n463_ = ~new_n64_ & ~new_n462_ & ~pi05;
  assign new_n464_ = ~pi10 & ~new_n62_ & ~pi09;
  assign new_n465_ = ~new_n463_ | ~new_n464_ | ~new_n37_ | ~pi14;
  assign new_n466_ = ~new_n24_ | ~pi02;
  assign new_n467_ = ~pi06 & ~pi05 & ~pi03 & ~new_n466_;
  assign new_n468_ = ~pi10 & ~new_n62_ & ~pi09;
  assign new_n469_ = ~new_n467_ | ~new_n468_ | ~new_n37_ | ~pi14;
  assign new_n470_ = ~pi02 | ~pi00;
  assign new_n471_ = ~pi06 & ~pi05 & ~pi03 & ~new_n470_;
  assign new_n472_ = ~pi10 & ~new_n62_ & ~pi09;
  assign new_n473_ = ~new_n471_ | ~new_n472_ | ~new_n37_ | ~pi14;
  assign new_n474_ = ~new_n461_ | ~new_n465_ | ~new_n469_ | ~new_n473_;
  assign new_n475_ = ~pi09 & ~pi10 & ~pi07;
  assign new_n476_ = ~new_n475_ | ~new_n37_ | ~pi14 | ~pi12;
  assign new_n477_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n478_ = ~new_n24_ | ~pi02;
  assign new_n479_ = ~new_n478_ & ~pi03 & ~new_n476_ & ~new_n477_;
  assign new_n480_ = ~pi09 & ~pi10;
  assign new_n481_ = ~pi12 | ~new_n480_ | ~new_n37_ | ~pi14;
  assign new_n482_ = ~pi02 | ~new_n66_ | ~new_n24_;
  assign new_n483_ = ~new_n56_ & ~pi06 & ~new_n481_ & ~new_n482_;
  assign new_n484_ = ~pi09 & ~pi10;
  assign new_n485_ = ~pi12 | ~new_n484_ | ~new_n37_ | ~pi14;
  assign new_n486_ = ~pi00 | ~new_n66_ | ~pi02;
  assign new_n487_ = ~new_n56_ & ~pi06 & ~new_n485_ & ~new_n486_;
  assign new_n488_ = ~new_n487_ & ~new_n483_ & ~new_n474_ & ~new_n479_;
  assign new_n489_ = ~new_n41_ & ~pi03 & ~new_n25_;
  assign new_n490_ = ~pi04 | ~new_n489_ | ~pi07;
  assign new_n491_ = ~pi08 | ~pi12 | ~new_n19_;
  assign new_n492_ = ~new_n27_ & ~pi15 & ~new_n490_ & ~new_n491_;
  assign new_n493_ = ~pi09 & ~pi10;
  assign new_n494_ = ~pi12 | ~new_n493_ | ~new_n37_ | ~pi14;
  assign new_n495_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n496_ = ~new_n56_ & ~new_n64_ & ~new_n494_ & ~new_n495_;
  assign new_n497_ = ~pi09 & ~pi10 & ~pi07;
  assign new_n498_ = ~new_n497_ | ~new_n37_ | ~pi14 | ~pi12;
  assign new_n499_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n500_ = ~new_n41_ | ~pi01;
  assign new_n501_ = ~new_n500_ & ~pi02 & ~new_n498_ & ~new_n499_;
  assign new_n502_ = ~pi09 & ~pi10 & ~pi07;
  assign new_n503_ = ~new_n502_ | ~new_n37_ | ~pi14 | ~pi12;
  assign new_n504_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n505_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n506_ = ~new_n505_ & ~new_n503_ & ~new_n504_;
  assign new_n507_ = ~new_n506_ & ~new_n501_ & ~new_n492_ & ~new_n496_;
  assign new_n508_ = ~pi09 & ~pi10;
  assign new_n509_ = ~pi12 | ~new_n508_ | ~new_n37_ | ~pi14;
  assign new_n510_ = ~pi01 | ~new_n25_ | ~new_n41_;
  assign new_n511_ = ~pi06 & ~pi05 & ~new_n509_ & ~new_n510_;
  assign new_n512_ = ~pi09 & ~pi10;
  assign new_n513_ = ~pi12 | ~new_n512_ | ~new_n37_ | ~pi14;
  assign new_n514_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n515_ = ~pi06 & ~pi05 & ~new_n513_ & ~new_n514_;
  assign new_n516_ = ~pi09 & ~pi10;
  assign new_n517_ = ~pi12 | ~new_n516_ | ~new_n37_ | ~pi14;
  assign new_n518_ = ~pi01 | ~new_n25_ | ~new_n41_;
  assign new_n519_ = ~new_n56_ & ~pi06 & ~new_n517_ & ~new_n518_;
  assign new_n520_ = ~pi09 & ~pi10;
  assign new_n521_ = ~pi12 | ~new_n520_ | ~new_n37_ | ~pi14;
  assign new_n522_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n523_ = ~new_n56_ & ~pi06 & ~new_n521_ & ~new_n522_;
  assign new_n524_ = ~new_n523_ & ~new_n519_ & ~new_n511_ & ~new_n515_;
  assign new_n525_ = ~new_n457_ | ~new_n488_ | ~new_n507_ | ~new_n524_;
  assign new_n526_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n527_ = ~pi06 & ~new_n526_ & ~pi05;
  assign new_n528_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n529_ = ~new_n527_ | ~new_n528_ | ~new_n27_ | ~pi13;
  assign new_n530_ = ~new_n57_ | ~pi04;
  assign new_n531_ = ~new_n24_ & ~pi00 & ~new_n530_ & ~pi02;
  assign new_n532_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n533_ = ~new_n531_ | ~new_n532_ | ~new_n27_ | ~pi13;
  assign new_n534_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n535_ = ~new_n56_ & ~new_n534_ & ~pi06;
  assign new_n536_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n537_ = ~new_n535_ | ~new_n536_ | ~new_n27_ | ~pi13;
  assign new_n538_ = ~new_n104_ | ~pi07;
  assign new_n539_ = ~new_n24_ & ~pi00 & ~new_n538_ & ~pi02;
  assign new_n540_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n541_ = ~new_n539_ | ~new_n540_ | ~new_n27_ | ~pi13;
  assign new_n542_ = ~new_n529_ | ~new_n533_ | ~new_n537_ | ~new_n541_;
  assign new_n543_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n544_ = ~new_n64_ & ~new_n543_ & ~pi05;
  assign new_n545_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n546_ = ~new_n544_ | ~new_n545_ | ~new_n27_ | ~pi13;
  assign new_n547_ = ~new_n24_ | ~pi02;
  assign new_n548_ = ~pi06 & ~pi05 & ~pi03 & ~new_n547_;
  assign new_n549_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n550_ = ~new_n548_ | ~new_n549_ | ~new_n27_ | ~pi13;
  assign new_n551_ = ~pi02 | ~pi00;
  assign new_n552_ = ~pi06 & ~pi05 & ~pi03 & ~new_n551_;
  assign new_n553_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n554_ = ~new_n552_ | ~new_n553_ | ~new_n27_ | ~pi13;
  assign new_n555_ = ~new_n57_ | ~pi04;
  assign new_n556_ = ~new_n25_ & ~pi01 & ~new_n555_ & ~pi03;
  assign new_n557_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n558_ = ~new_n556_ | ~new_n557_ | ~new_n27_ | ~pi13;
  assign new_n559_ = ~new_n546_ | ~new_n550_ | ~new_n554_ | ~new_n558_;
  assign new_n560_ = ~pi02 | ~pi00;
  assign new_n561_ = ~new_n56_ & ~pi06 & ~pi03 & ~new_n560_;
  assign new_n562_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n563_ = ~new_n561_ | ~new_n562_ | ~new_n27_ | ~pi13;
  assign new_n564_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n565_ = ~new_n25_ & ~pi01 & ~new_n564_ & ~pi03;
  assign new_n566_ = ~pi09 & ~pi10 & ~pi07;
  assign new_n567_ = ~new_n26_ & ~pi14 & ~pi12;
  assign new_n568_ = ~new_n567_ | ~new_n565_ | ~new_n566_;
  assign new_n569_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n570_ = ~new_n41_ & ~new_n25_ & ~new_n569_ & ~pi03;
  assign new_n571_ = ~pi09 & ~pi10 & ~pi07;
  assign new_n572_ = ~new_n26_ & ~pi14 & ~pi12;
  assign new_n573_ = ~new_n572_ | ~new_n570_ | ~new_n571_;
  assign new_n574_ = ~new_n104_ | ~pi07;
  assign new_n575_ = ~new_n25_ & ~pi01 & ~new_n574_ & ~pi03;
  assign new_n576_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n577_ = ~new_n575_ | ~new_n576_ | ~new_n27_ | ~pi13;
  assign new_n578_ = ~new_n563_ | ~new_n568_ | ~new_n573_ | ~new_n577_;
  assign new_n579_ = ~pi07 | ~pi04;
  assign new_n580_ = ~new_n41_ & ~new_n25_ & ~new_n579_ & ~pi03;
  assign new_n581_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n582_ = ~new_n580_ | ~new_n581_ | ~new_n27_ | ~pi13;
  assign new_n583_ = ~pi02 | ~pi00;
  assign new_n584_ = ~new_n64_ & ~pi05 & ~pi03 & ~new_n583_;
  assign new_n585_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n586_ = ~new_n584_ | ~new_n585_ | ~new_n27_ | ~pi13;
  assign new_n587_ = ~pi07 | ~pi04;
  assign new_n588_ = ~new_n25_ & ~pi01 & ~new_n587_ & ~pi03;
  assign new_n589_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n590_ = ~new_n588_ | ~new_n589_ | ~new_n27_ | ~pi13;
  assign new_n591_ = ~new_n590_ | ~new_n582_ | ~new_n586_;
  assign new_n592_ = ~new_n591_ & ~new_n578_ & ~new_n542_ & ~new_n559_;
  assign new_n593_ = ~pi07 | ~pi04;
  assign new_n594_ = ~new_n24_ & ~pi00 & ~new_n593_ & ~pi02;
  assign new_n595_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n596_ = ~new_n594_ | ~new_n595_ | ~new_n27_ | ~pi13;
  assign new_n597_ = ~pi07 | ~pi04;
  assign new_n598_ = ~new_n25_ & ~pi01 & ~new_n597_ & ~pi03;
  assign new_n599_ = ~pi10 & ~pi13 & ~pi09;
  assign new_n600_ = ~new_n598_ | ~new_n599_ | ~new_n37_ | ~pi14;
  assign new_n601_ = ~pi07 | ~pi04;
  assign new_n602_ = ~new_n41_ & ~new_n25_ & ~new_n601_ & ~pi03;
  assign new_n603_ = ~pi10 & ~pi13 & ~pi09;
  assign new_n604_ = ~new_n602_ | ~new_n603_ | ~new_n37_ | ~pi14;
  assign new_n605_ = ~pi07 | ~pi04;
  assign new_n606_ = ~new_n24_ & ~pi00 & ~new_n605_ & ~new_n66_;
  assign new_n607_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n608_ = ~new_n606_ | ~new_n607_ | ~new_n27_ | ~pi13;
  assign new_n609_ = ~new_n596_ | ~new_n600_ | ~new_n604_ | ~new_n608_;
  assign new_n610_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n611_ = ~pi13 | ~new_n610_ | ~new_n27_;
  assign new_n612_ = ~pi01 | ~new_n25_ | ~new_n41_;
  assign new_n613_ = ~pi06 & ~pi05 & ~new_n611_ & ~new_n612_;
  assign new_n614_ = ~pi09 & ~pi10 & ~pi07;
  assign new_n615_ = ~new_n614_ | ~new_n27_ | ~new_n62_ | ~pi13;
  assign new_n616_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n617_ = ~new_n41_ | ~pi01;
  assign new_n618_ = ~new_n617_ & ~pi02 & ~new_n615_ & ~new_n616_;
  assign new_n619_ = ~pi09 & ~pi10 & ~pi07;
  assign new_n620_ = ~new_n619_ | ~new_n27_ | ~new_n62_ | ~pi13;
  assign new_n621_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n622_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n623_ = ~new_n622_ & ~new_n620_ & ~new_n621_;
  assign new_n624_ = ~new_n623_ & ~new_n618_ & ~new_n609_ & ~new_n613_;
  assign new_n625_ = ~pi10 & ~pi13 & ~pi09;
  assign new_n626_ = ~pi14 | ~new_n625_ | ~new_n37_;
  assign new_n627_ = ~pi02 | ~new_n66_ | ~new_n24_;
  assign new_n628_ = ~pi06 & ~pi05 & ~new_n626_ & ~new_n627_;
  assign new_n629_ = ~pi10 & ~pi13 & ~pi09;
  assign new_n630_ = ~pi14 | ~new_n629_ | ~new_n37_;
  assign new_n631_ = ~pi00 | ~new_n66_ | ~pi02;
  assign new_n632_ = ~pi06 & ~pi05 & ~new_n630_ & ~new_n631_;
  assign new_n633_ = ~pi10 & ~pi13 & ~pi09;
  assign new_n634_ = ~pi14 | ~new_n633_ | ~new_n37_;
  assign new_n635_ = ~pi02 | ~new_n66_ | ~new_n24_;
  assign new_n636_ = ~new_n56_ & ~pi06 & ~new_n634_ & ~new_n635_;
  assign new_n637_ = ~pi10 & ~pi13 & ~pi09;
  assign new_n638_ = ~pi14 | ~new_n637_ | ~new_n37_;
  assign new_n639_ = ~pi00 | ~new_n66_ | ~pi02;
  assign new_n640_ = ~new_n56_ & ~pi06 & ~new_n638_ & ~new_n639_;
  assign new_n641_ = ~new_n640_ & ~new_n636_ & ~new_n628_ & ~new_n632_;
  assign new_n642_ = ~pi09 & ~pi10 & ~pi07;
  assign new_n643_ = ~new_n642_ | ~new_n37_ | ~new_n26_ | ~pi14;
  assign new_n644_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n645_ = ~new_n24_ | ~pi02;
  assign new_n646_ = ~new_n645_ & ~pi03 & ~new_n643_ & ~new_n644_;
  assign new_n647_ = ~pi09 & ~pi10 & ~pi07;
  assign new_n648_ = ~new_n647_ | ~new_n37_ | ~new_n26_ | ~pi14;
  assign new_n649_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n650_ = ~pi02 | ~pi00;
  assign new_n651_ = ~new_n650_ & ~pi03 & ~new_n648_ & ~new_n649_;
  assign new_n652_ = ~pi10 & ~pi13 & ~pi09;
  assign new_n653_ = ~pi14 | ~new_n652_ | ~new_n37_;
  assign new_n654_ = ~pi02 | ~new_n66_ | ~new_n24_;
  assign new_n655_ = ~new_n64_ & ~pi05 & ~new_n653_ & ~new_n654_;
  assign new_n656_ = ~pi10 & ~pi13 & ~pi09;
  assign new_n657_ = ~pi14 | ~new_n656_ | ~new_n37_;
  assign new_n658_ = ~pi00 | ~new_n66_ | ~pi02;
  assign new_n659_ = ~new_n64_ & ~pi05 & ~new_n657_ & ~new_n658_;
  assign new_n660_ = ~new_n659_ & ~new_n655_ & ~new_n646_ & ~new_n651_;
  assign new_n661_ = ~new_n592_ | ~new_n624_ | ~new_n641_ | ~new_n660_;
  assign new_n662_ = ~new_n27_ & ~pi15 & ~pi13;
  assign new_n663_ = ~new_n662_ | ~pi11 | ~new_n64_ | ~pi08;
  assign new_n664_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n665_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n666_ = ~new_n665_ & ~new_n663_ & ~new_n664_;
  assign new_n667_ = ~pi05 & ~pi06;
  assign new_n668_ = ~new_n667_ | ~new_n25_ | ~new_n41_ | ~pi01;
  assign new_n669_ = ~pi11 | ~new_n26_ | ~pi08;
  assign new_n670_ = ~new_n27_ & ~pi15 & ~new_n668_ & ~new_n669_;
  assign new_n671_ = ~pi05 & ~pi06;
  assign new_n672_ = ~new_n671_ | ~pi03 | ~new_n41_ | ~pi01;
  assign new_n673_ = ~pi11 | ~new_n26_ | ~pi08;
  assign new_n674_ = ~new_n27_ & ~pi15 & ~new_n672_ & ~new_n673_;
  assign new_n675_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n676_ = ~pi04 | ~new_n675_ | ~new_n57_;
  assign new_n677_ = ~pi11 | ~new_n26_ | ~pi08;
  assign new_n678_ = ~new_n27_ & ~pi15 & ~new_n676_ & ~new_n677_;
  assign new_n679_ = ~new_n678_ & ~new_n674_ & ~new_n666_ & ~new_n670_;
  assign new_n680_ = ~pi08 | ~pi11;
  assign new_n681_ = ~new_n27_ & ~pi15 & ~pi13 & ~new_n680_;
  assign new_n682_ = ~new_n24_ & ~new_n66_ & ~pi00;
  assign new_n683_ = ~new_n681_ | ~new_n682_ | ~new_n104_ | ~pi07;
  assign new_n684_ = ~pi08 | ~pi11;
  assign new_n685_ = ~new_n27_ & ~pi15 & ~pi13 & ~new_n684_;
  assign new_n686_ = ~new_n24_ & ~new_n66_ & ~pi00;
  assign new_n687_ = ~new_n685_ | ~new_n686_ | ~new_n57_ | ~pi04;
  assign new_n688_ = ~pi08 | ~pi11;
  assign new_n689_ = ~new_n27_ & ~pi15 & ~pi13 & ~new_n688_;
  assign new_n690_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n691_ = ~new_n689_ | ~new_n690_ | ~new_n104_ | ~pi07;
  assign new_n692_ = ~new_n679_ | ~new_n683_ | ~new_n687_ | ~new_n691_;
  assign new_n693_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n694_ = ~new_n41_ & ~new_n25_ & ~new_n693_ & ~pi03;
  assign new_n695_ = ~new_n62_ & ~pi15 & ~new_n27_;
  assign new_n696_ = ~pi07 & ~pi09;
  assign new_n697_ = ~new_n694_ | ~new_n695_ | ~pi11 | ~new_n696_;
  assign new_n698_ = ~pi11 | ~pi12 | ~new_n79_;
  assign new_n699_ = ~new_n27_ & ~new_n698_ & ~pi15;
  assign new_n700_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n701_ = ~new_n699_ | ~new_n700_ | ~new_n104_ | ~pi07;
  assign new_n702_ = ~pi02 | ~pi00;
  assign new_n703_ = ~new_n64_ & ~pi05 & ~pi03 & ~new_n702_;
  assign new_n704_ = ~new_n22_ & ~new_n62_ & ~pi09;
  assign new_n705_ = ~new_n703_ | ~new_n704_ | ~new_n37_ | ~pi14;
  assign new_n706_ = ~pi11 | ~pi12 | ~new_n79_;
  assign new_n707_ = ~new_n27_ & ~new_n706_ & ~pi15;
  assign new_n708_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n709_ = ~new_n707_ | ~new_n708_ | ~pi07 | ~pi04;
  assign new_n710_ = ~new_n697_ | ~new_n701_ | ~new_n705_ | ~new_n709_;
  assign new_n711_ = ~pi11 | ~pi12 | ~new_n79_;
  assign new_n712_ = ~new_n27_ & ~new_n711_ & ~pi15;
  assign new_n713_ = ~new_n41_ & ~pi03 & ~new_n25_;
  assign new_n714_ = ~new_n712_ | ~new_n713_ | ~pi07 | ~pi04;
  assign new_n715_ = ~pi08 | ~pi11;
  assign new_n716_ = ~new_n27_ & ~pi15 & ~pi13 & ~new_n715_;
  assign new_n717_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n718_ = ~new_n716_ | ~new_n717_ | ~pi07 | ~pi04;
  assign new_n719_ = ~pi08 | ~pi11;
  assign new_n720_ = ~new_n27_ & ~pi15 & ~pi13 & ~new_n719_;
  assign new_n721_ = ~new_n24_ & ~new_n66_ & ~pi00;
  assign new_n722_ = ~new_n720_ | ~new_n721_ | ~pi07 | ~pi04;
  assign new_n723_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n724_ = ~new_n24_ & ~pi00 & ~new_n723_ & ~pi02;
  assign new_n725_ = ~pi08 | ~pi11 | ~new_n64_;
  assign new_n726_ = ~new_n27_ & ~pi13 & ~new_n725_ & ~pi15;
  assign new_n727_ = ~new_n724_ | ~new_n726_;
  assign new_n728_ = ~new_n714_ | ~new_n718_ | ~new_n722_ | ~new_n727_;
  assign new_n729_ = ~new_n728_ & ~new_n692_ & ~new_n710_;
  assign new_n730_ = ~pi11 | ~pi12 | ~new_n79_;
  assign new_n731_ = ~new_n27_ & ~new_n730_ & ~pi15;
  assign new_n732_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n733_ = ~new_n731_ | ~new_n732_ | ~new_n104_ | ~pi07;
  assign new_n734_ = ~pi11 | ~pi12 | ~new_n79_;
  assign new_n735_ = ~new_n27_ & ~new_n734_ & ~pi15;
  assign new_n736_ = ~new_n24_ & ~new_n66_ & ~pi00;
  assign new_n737_ = ~new_n735_ | ~new_n736_ | ~new_n104_ | ~pi07;
  assign new_n738_ = ~new_n24_ | ~pi02;
  assign new_n739_ = ~pi06 & ~pi05 & ~pi03 & ~new_n738_;
  assign new_n740_ = ~new_n22_ & ~new_n62_ & ~pi09;
  assign new_n741_ = ~new_n739_ | ~new_n740_ | ~new_n37_ | ~pi14;
  assign new_n742_ = ~pi02 | ~pi00;
  assign new_n743_ = ~pi06 & ~pi05 & ~pi03 & ~new_n742_;
  assign new_n744_ = ~new_n22_ & ~new_n62_ & ~pi09;
  assign new_n745_ = ~new_n743_ | ~new_n744_ | ~new_n37_ | ~pi14;
  assign new_n746_ = ~new_n733_ | ~new_n737_ | ~new_n741_ | ~new_n745_;
  assign new_n747_ = ~pi09 & ~new_n22_ & ~pi07;
  assign new_n748_ = ~new_n747_ | ~new_n37_ | ~pi14 | ~pi12;
  assign new_n749_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n750_ = ~new_n24_ | ~pi02;
  assign new_n751_ = ~new_n750_ & ~pi03 & ~new_n748_ & ~new_n749_;
  assign new_n752_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n753_ = ~pi04 | ~new_n752_ | ~new_n57_;
  assign new_n754_ = ~pi11 | ~pi12 | ~new_n79_;
  assign new_n755_ = ~new_n27_ & ~pi15 & ~new_n753_ & ~new_n754_;
  assign new_n756_ = ~pi06 & ~new_n56_;
  assign new_n757_ = ~new_n756_ | ~new_n66_ | ~pi02 | ~pi00;
  assign new_n758_ = ~pi11 | ~pi12 | ~new_n79_;
  assign new_n759_ = ~new_n27_ & ~pi15 & ~new_n757_ & ~new_n758_;
  assign new_n760_ = ~new_n759_ & ~new_n755_ & ~new_n746_ & ~new_n751_;
  assign new_n761_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n762_ = ~pi04 | ~new_n761_ | ~pi07;
  assign new_n763_ = ~pi11 | ~pi12 | ~new_n79_;
  assign new_n764_ = ~new_n27_ & ~pi15 & ~new_n762_ & ~new_n763_;
  assign new_n765_ = ~pi00 & ~new_n24_;
  assign new_n766_ = ~pi03 | ~new_n765_ | ~pi07 | ~pi04;
  assign new_n767_ = ~pi11 | ~pi12 | ~new_n79_;
  assign new_n768_ = ~new_n27_ & ~pi15 & ~new_n766_ & ~new_n767_;
  assign new_n769_ = ~pi09 & ~new_n22_ & ~pi07;
  assign new_n770_ = ~new_n769_ | ~new_n37_ | ~pi14 | ~pi12;
  assign new_n771_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n772_ = ~new_n41_ | ~pi01;
  assign new_n773_ = ~new_n772_ & ~pi02 & ~new_n770_ & ~new_n771_;
  assign new_n774_ = ~pi09 & ~new_n22_ & ~pi07;
  assign new_n775_ = ~new_n774_ | ~new_n37_ | ~pi14 | ~pi12;
  assign new_n776_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n777_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n778_ = ~new_n777_ & ~new_n775_ & ~new_n776_;
  assign new_n779_ = ~new_n778_ & ~new_n773_ & ~new_n764_ & ~new_n768_;
  assign new_n780_ = ~pi05 & ~pi06;
  assign new_n781_ = ~new_n780_ | ~new_n25_ | ~new_n41_ | ~pi01;
  assign new_n782_ = ~pi11 | ~pi12 | ~new_n79_;
  assign new_n783_ = ~new_n27_ & ~pi15 & ~new_n781_ & ~new_n782_;
  assign new_n784_ = ~pi05 & ~pi06;
  assign new_n785_ = ~new_n784_ | ~pi03 | ~new_n41_ | ~pi01;
  assign new_n786_ = ~pi11 | ~pi12 | ~new_n79_;
  assign new_n787_ = ~new_n27_ & ~pi15 & ~new_n785_ & ~new_n786_;
  assign new_n788_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n789_ = ~pi04 | ~new_n788_ | ~new_n57_;
  assign new_n790_ = ~pi11 | ~pi12 | ~new_n79_;
  assign new_n791_ = ~new_n27_ & ~pi15 & ~new_n789_ & ~new_n790_;
  assign new_n792_ = ~pi06 & ~new_n56_;
  assign new_n793_ = ~new_n792_ | ~pi03 | ~new_n41_ | ~pi01;
  assign new_n794_ = ~pi11 | ~pi12 | ~new_n79_;
  assign new_n795_ = ~new_n27_ & ~pi15 & ~new_n793_ & ~new_n794_;
  assign new_n796_ = ~new_n795_ & ~new_n791_ & ~new_n783_ & ~new_n787_;
  assign new_n797_ = ~new_n729_ | ~new_n760_ | ~new_n779_ | ~new_n796_;
  assign new_n798_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n799_ = ~pi06 & ~new_n798_ & ~pi05;
  assign new_n800_ = ~new_n89_ & ~pi13 & ~pi10;
  assign new_n801_ = ~new_n799_ | ~new_n800_ | ~new_n37_ | ~pi14;
  assign new_n802_ = ~new_n57_ | ~pi04;
  assign new_n803_ = ~new_n24_ & ~pi00 & ~new_n802_ & ~pi02;
  assign new_n804_ = ~new_n89_ & ~pi13 & ~pi10;
  assign new_n805_ = ~new_n803_ | ~new_n804_ | ~new_n37_ | ~pi14;
  assign new_n806_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n807_ = ~new_n56_ & ~new_n806_ & ~pi06;
  assign new_n808_ = ~new_n89_ & ~pi13 & ~pi10;
  assign new_n809_ = ~new_n807_ | ~new_n808_ | ~new_n37_ | ~pi14;
  assign new_n810_ = ~new_n104_ | ~pi07;
  assign new_n811_ = ~new_n24_ & ~pi00 & ~new_n810_ & ~pi02;
  assign new_n812_ = ~new_n89_ & ~pi13 & ~pi10;
  assign new_n813_ = ~new_n811_ | ~new_n812_ | ~new_n37_ | ~pi14;
  assign new_n814_ = ~new_n801_ | ~new_n805_ | ~new_n809_ | ~new_n813_;
  assign new_n815_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n816_ = ~new_n64_ & ~new_n815_ & ~pi05;
  assign new_n817_ = ~new_n89_ & ~pi13 & ~pi10;
  assign new_n818_ = ~new_n816_ | ~new_n817_ | ~new_n37_ | ~pi14;
  assign new_n819_ = ~new_n24_ | ~pi02;
  assign new_n820_ = ~pi06 & ~pi05 & ~pi03 & ~new_n819_;
  assign new_n821_ = ~new_n89_ & ~pi13 & ~pi10;
  assign new_n822_ = ~new_n820_ | ~new_n821_ | ~new_n37_ | ~pi14;
  assign new_n823_ = ~pi02 | ~pi00;
  assign new_n824_ = ~pi06 & ~pi05 & ~pi03 & ~new_n823_;
  assign new_n825_ = ~new_n89_ & ~pi13 & ~pi10;
  assign new_n826_ = ~new_n824_ | ~new_n825_ | ~new_n37_ | ~pi14;
  assign new_n827_ = ~new_n57_ | ~pi04;
  assign new_n828_ = ~new_n25_ & ~pi01 & ~new_n827_ & ~pi03;
  assign new_n829_ = ~new_n89_ & ~pi13 & ~pi10;
  assign new_n830_ = ~new_n828_ | ~new_n829_ | ~new_n37_ | ~pi14;
  assign new_n831_ = ~new_n818_ | ~new_n822_ | ~new_n826_ | ~new_n830_;
  assign new_n832_ = ~pi02 | ~pi00;
  assign new_n833_ = ~new_n56_ & ~pi06 & ~pi03 & ~new_n832_;
  assign new_n834_ = ~new_n89_ & ~pi13 & ~pi10;
  assign new_n835_ = ~new_n833_ | ~new_n834_ | ~new_n37_ | ~pi14;
  assign new_n836_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n837_ = ~new_n25_ & ~pi01 & ~new_n836_ & ~pi03;
  assign new_n838_ = ~new_n89_ & ~pi10 & ~pi07;
  assign new_n839_ = ~new_n27_ & ~pi15 & ~pi13;
  assign new_n840_ = ~new_n839_ | ~new_n837_ | ~new_n838_;
  assign new_n841_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n842_ = ~new_n41_ & ~new_n25_ & ~new_n841_ & ~pi03;
  assign new_n843_ = ~new_n89_ & ~pi10 & ~pi07;
  assign new_n844_ = ~new_n27_ & ~pi15 & ~pi13;
  assign new_n845_ = ~new_n844_ | ~new_n842_ | ~new_n843_;
  assign new_n846_ = ~new_n104_ | ~pi07;
  assign new_n847_ = ~new_n25_ & ~pi01 & ~new_n846_ & ~pi03;
  assign new_n848_ = ~new_n89_ & ~pi13 & ~pi10;
  assign new_n849_ = ~new_n847_ | ~new_n848_ | ~new_n37_ | ~pi14;
  assign new_n850_ = ~new_n835_ | ~new_n840_ | ~new_n845_ | ~new_n849_;
  assign new_n851_ = ~pi07 | ~pi04;
  assign new_n852_ = ~new_n41_ & ~new_n25_ & ~new_n851_ & ~pi03;
  assign new_n853_ = ~new_n89_ & ~pi13 & ~pi10;
  assign new_n854_ = ~new_n852_ | ~new_n853_ | ~new_n37_ | ~pi14;
  assign new_n855_ = ~pi02 | ~pi00;
  assign new_n856_ = ~new_n64_ & ~pi05 & ~pi03 & ~new_n855_;
  assign new_n857_ = ~new_n89_ & ~pi13 & ~pi10;
  assign new_n858_ = ~new_n856_ | ~new_n857_ | ~new_n37_ | ~pi14;
  assign new_n859_ = ~pi07 | ~pi04;
  assign new_n860_ = ~new_n25_ & ~pi01 & ~new_n859_ & ~pi03;
  assign new_n861_ = ~new_n89_ & ~pi13 & ~pi10;
  assign new_n862_ = ~new_n860_ | ~new_n861_ | ~new_n37_ | ~pi14;
  assign new_n863_ = ~new_n862_ | ~new_n854_ | ~new_n858_;
  assign new_n864_ = ~new_n863_ & ~new_n850_ & ~new_n814_ & ~new_n831_;
  assign new_n865_ = ~pi07 | ~pi04;
  assign new_n866_ = ~new_n24_ & ~pi00 & ~new_n865_ & ~pi02;
  assign new_n867_ = ~new_n89_ & ~pi13 & ~pi10;
  assign new_n868_ = ~new_n866_ | ~new_n867_ | ~new_n37_ | ~pi14;
  assign new_n869_ = ~pi08 | ~pi11;
  assign new_n870_ = ~new_n27_ & ~pi15 & ~pi13 & ~new_n869_;
  assign new_n871_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n872_ = ~new_n870_ | ~new_n871_ | ~pi07 | ~pi04;
  assign new_n873_ = ~pi08 | ~pi11;
  assign new_n874_ = ~new_n27_ & ~pi15 & ~pi13 & ~new_n873_;
  assign new_n875_ = ~new_n41_ & ~pi03 & ~new_n25_;
  assign new_n876_ = ~new_n874_ | ~new_n875_ | ~pi07 | ~pi04;
  assign new_n877_ = ~pi07 | ~pi04;
  assign new_n878_ = ~new_n24_ & ~pi00 & ~new_n877_ & ~new_n66_;
  assign new_n879_ = ~new_n89_ & ~pi13 & ~pi10;
  assign new_n880_ = ~new_n878_ | ~new_n879_ | ~new_n37_ | ~pi14;
  assign new_n881_ = ~new_n868_ | ~new_n872_ | ~new_n876_ | ~new_n880_;
  assign new_n882_ = ~new_n89_ & ~pi13 & ~pi10;
  assign new_n883_ = ~pi14 | ~new_n882_ | ~new_n37_;
  assign new_n884_ = ~pi01 | ~new_n25_ | ~new_n41_;
  assign new_n885_ = ~pi06 & ~pi05 & ~new_n883_ & ~new_n884_;
  assign new_n886_ = ~new_n89_ & ~pi10 & ~pi07;
  assign new_n887_ = ~new_n886_ | ~new_n37_ | ~new_n26_ | ~pi14;
  assign new_n888_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n889_ = ~new_n41_ | ~pi01;
  assign new_n890_ = ~new_n889_ & ~pi02 & ~new_n887_ & ~new_n888_;
  assign new_n891_ = ~new_n89_ & ~pi10 & ~pi07;
  assign new_n892_ = ~new_n891_ | ~new_n37_ | ~new_n26_ | ~pi14;
  assign new_n893_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n894_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n895_ = ~new_n894_ & ~new_n892_ & ~new_n893_;
  assign new_n896_ = ~new_n895_ & ~new_n890_ & ~new_n881_ & ~new_n885_;
  assign new_n897_ = ~pi05 & ~pi06;
  assign new_n898_ = ~new_n897_ | ~new_n66_ | ~new_n24_ | ~pi02;
  assign new_n899_ = ~pi11 | ~new_n26_ | ~pi08;
  assign new_n900_ = ~new_n27_ & ~pi15 & ~new_n898_ & ~new_n899_;
  assign new_n901_ = ~pi05 & ~pi06;
  assign new_n902_ = ~new_n901_ | ~new_n66_ | ~pi02 | ~pi00;
  assign new_n903_ = ~pi11 | ~new_n26_ | ~pi08;
  assign new_n904_ = ~new_n27_ & ~pi15 & ~new_n902_ & ~new_n903_;
  assign new_n905_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n906_ = ~pi04 | ~new_n905_ | ~new_n57_;
  assign new_n907_ = ~pi11 | ~new_n26_ | ~pi08;
  assign new_n908_ = ~new_n27_ & ~pi15 & ~new_n906_ & ~new_n907_;
  assign new_n909_ = ~pi06 & ~new_n56_;
  assign new_n910_ = ~new_n909_ | ~new_n66_ | ~pi02 | ~pi00;
  assign new_n911_ = ~pi11 | ~new_n26_ | ~pi08;
  assign new_n912_ = ~new_n27_ & ~pi15 & ~new_n910_ & ~new_n911_;
  assign new_n913_ = ~new_n912_ & ~new_n908_ & ~new_n900_ & ~new_n904_;
  assign new_n914_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n915_ = ~new_n914_ | ~pi06 | ~new_n56_ | ~pi05;
  assign new_n916_ = ~new_n27_ & ~pi15 & ~pi13;
  assign new_n917_ = ~new_n916_ | ~pi11 | ~new_n64_ | ~pi08;
  assign new_n918_ = ~new_n915_ & ~new_n917_;
  assign new_n919_ = ~new_n27_ & ~pi15 & ~pi13;
  assign new_n920_ = ~new_n919_ | ~pi11 | ~new_n64_ | ~pi08;
  assign new_n921_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n922_ = ~pi02 | ~pi00;
  assign new_n923_ = ~new_n922_ & ~pi03 & ~new_n920_ & ~new_n921_;
  assign new_n924_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n925_ = ~pi07 | ~new_n924_ | ~new_n104_;
  assign new_n926_ = ~pi11 | ~new_n26_ | ~pi08;
  assign new_n927_ = ~new_n27_ & ~pi15 & ~new_n925_ & ~new_n926_;
  assign new_n928_ = ~pi05 & ~new_n64_;
  assign new_n929_ = ~new_n928_ | ~new_n66_ | ~pi02 | ~pi00;
  assign new_n930_ = ~pi11 | ~new_n26_ | ~pi08;
  assign new_n931_ = ~new_n27_ & ~pi15 & ~new_n929_ & ~new_n930_;
  assign new_n932_ = ~new_n931_ & ~new_n927_ & ~new_n918_ & ~new_n923_;
  assign new_n933_ = ~new_n864_ | ~new_n896_ | ~new_n913_ | ~new_n932_;
  assign new_n934_ = ~new_n933_ & ~new_n797_ & ~new_n525_ & ~new_n661_;
  assign new_n935_ = ~pi07 | ~pi04;
  assign new_n936_ = ~new_n24_ & ~pi00 & ~new_n935_ & ~pi02;
  assign new_n937_ = ~new_n22_ & ~pi13 & ~pi09;
  assign new_n938_ = ~new_n936_ | ~new_n937_ | ~new_n37_ | ~pi14;
  assign new_n939_ = ~pi07 | ~pi04;
  assign new_n940_ = ~new_n24_ & ~pi00 & ~new_n939_ & ~new_n66_;
  assign new_n941_ = ~new_n22_ & ~pi13 & ~pi09;
  assign new_n942_ = ~new_n940_ | ~new_n941_ | ~new_n37_ | ~pi14;
  assign new_n943_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n944_ = ~new_n24_ & ~pi00 & ~new_n943_ & ~pi02;
  assign new_n945_ = ~new_n27_ & ~pi15 & ~pi13;
  assign new_n946_ = ~pi07 & ~pi09;
  assign new_n947_ = ~new_n944_ | ~new_n945_ | ~pi11 | ~new_n946_;
  assign new_n948_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n949_ = ~new_n24_ & ~pi00 & ~new_n948_ & ~new_n66_;
  assign new_n950_ = ~new_n27_ & ~pi15 & ~pi13;
  assign new_n951_ = ~pi07 & ~pi09;
  assign new_n952_ = ~new_n949_ | ~new_n950_ | ~pi11 | ~new_n951_;
  assign new_n953_ = ~new_n938_ | ~new_n942_ | ~new_n947_ | ~new_n952_;
  assign new_n954_ = ~new_n41_ | ~pi01;
  assign new_n955_ = ~pi06 & ~pi05 & ~pi02 & ~new_n954_;
  assign new_n956_ = ~new_n22_ & ~pi13 & ~pi09;
  assign new_n957_ = ~new_n955_ | ~new_n956_ | ~new_n37_ | ~pi14;
  assign new_n958_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n959_ = ~pi06 & ~new_n958_ & ~pi05;
  assign new_n960_ = ~new_n22_ & ~pi13 & ~pi09;
  assign new_n961_ = ~new_n959_ | ~new_n960_ | ~new_n37_ | ~pi14;
  assign new_n962_ = ~new_n57_ | ~pi04;
  assign new_n963_ = ~new_n24_ & ~pi00 & ~new_n962_ & ~pi02;
  assign new_n964_ = ~new_n22_ & ~pi13 & ~pi09;
  assign new_n965_ = ~new_n963_ | ~new_n964_ | ~new_n37_ | ~pi14;
  assign new_n966_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n967_ = ~new_n56_ & ~new_n966_ & ~pi06;
  assign new_n968_ = ~new_n22_ & ~pi13 & ~pi09;
  assign new_n969_ = ~new_n967_ | ~new_n968_ | ~new_n37_ | ~pi14;
  assign new_n970_ = ~new_n957_ | ~new_n961_ | ~new_n965_ | ~new_n969_;
  assign new_n971_ = ~new_n104_ | ~pi07;
  assign new_n972_ = ~new_n24_ & ~pi00 & ~new_n971_ & ~pi02;
  assign new_n973_ = ~new_n22_ & ~pi13 & ~pi09;
  assign new_n974_ = ~new_n972_ | ~new_n973_ | ~new_n37_ | ~pi14;
  assign new_n975_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n976_ = ~new_n64_ & ~new_n975_ & ~pi05;
  assign new_n977_ = ~new_n22_ & ~pi13 & ~pi09;
  assign new_n978_ = ~new_n976_ | ~new_n977_ | ~new_n37_ | ~pi14;
  assign new_n979_ = ~new_n24_ | ~pi02;
  assign new_n980_ = ~pi06 & ~pi05 & ~pi03 & ~new_n979_;
  assign new_n981_ = ~new_n22_ & ~pi13 & ~pi09;
  assign new_n982_ = ~new_n980_ | ~new_n981_ | ~new_n37_ | ~pi14;
  assign new_n983_ = ~pi02 | ~pi00;
  assign new_n984_ = ~pi06 & ~pi05 & ~pi03 & ~new_n983_;
  assign new_n985_ = ~new_n22_ & ~pi13 & ~pi09;
  assign new_n986_ = ~new_n984_ | ~new_n985_ | ~new_n37_ | ~pi14;
  assign new_n987_ = ~new_n974_ | ~new_n978_ | ~new_n982_ | ~new_n986_;
  assign new_n988_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n989_ = ~new_n25_ & ~pi01 & ~new_n988_ & ~pi03;
  assign new_n990_ = ~new_n27_ & ~pi15 & ~pi13;
  assign new_n991_ = ~pi07 & ~pi09;
  assign new_n992_ = ~new_n989_ | ~new_n990_ | ~pi11 | ~new_n991_;
  assign new_n993_ = ~new_n57_ | ~pi04;
  assign new_n994_ = ~new_n25_ & ~pi01 & ~new_n993_ & ~pi03;
  assign new_n995_ = ~new_n22_ & ~pi13 & ~pi09;
  assign new_n996_ = ~new_n994_ | ~new_n995_ | ~new_n37_ | ~pi14;
  assign new_n997_ = ~pi02 | ~pi00;
  assign new_n998_ = ~new_n56_ & ~pi06 & ~pi03 & ~new_n997_;
  assign new_n999_ = ~new_n22_ & ~pi13 & ~pi09;
  assign new_n1000_ = ~new_n998_ | ~new_n999_ | ~new_n37_ | ~pi14;
  assign new_n1001_ = ~new_n1000_ | ~new_n992_ | ~new_n996_;
  assign new_n1002_ = ~new_n1001_ & ~new_n987_ & ~new_n953_ & ~new_n970_;
  assign new_n1003_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1004_ = ~new_n24_ & ~pi00 & ~new_n1003_ & ~new_n66_;
  assign new_n1005_ = ~new_n26_ & ~pi14 & ~pi12;
  assign new_n1006_ = ~pi07 & ~pi09;
  assign new_n1007_ = ~new_n1004_ | ~new_n1005_ | ~pi11 | ~new_n1006_;
  assign new_n1008_ = ~new_n41_ | ~pi01;
  assign new_n1009_ = ~pi06 & ~pi05 & ~pi02 & ~new_n1008_;
  assign new_n1010_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1011_ = ~new_n1009_ | ~new_n1010_ | ~new_n27_ | ~pi13;
  assign new_n1012_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1013_ = ~pi06 & ~new_n1012_ & ~pi05;
  assign new_n1014_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1015_ = ~new_n1013_ | ~new_n1014_ | ~new_n27_ | ~pi13;
  assign new_n1016_ = ~new_n57_ | ~pi04;
  assign new_n1017_ = ~new_n24_ & ~pi00 & ~new_n1016_ & ~pi02;
  assign new_n1018_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1019_ = ~new_n1017_ | ~new_n1018_ | ~new_n27_ | ~pi13;
  assign new_n1020_ = ~new_n1007_ | ~new_n1011_ | ~new_n1015_ | ~new_n1019_;
  assign new_n1021_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1022_ = ~pi13 | ~new_n1021_ | ~new_n27_;
  assign new_n1023_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1024_ = ~new_n64_ & ~pi05 & ~new_n1022_ & ~new_n1023_;
  assign new_n1025_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1026_ = ~pi13 | ~new_n1025_ | ~new_n27_;
  assign new_n1027_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1028_ = ~new_n56_ & ~pi06 & ~new_n1026_ & ~new_n1027_;
  assign new_n1029_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1030_ = ~pi13 | ~new_n1029_ | ~new_n27_;
  assign new_n1031_ = ~pi01 | ~new_n25_ | ~new_n41_;
  assign new_n1032_ = ~new_n64_ & ~pi05 & ~new_n1030_ & ~new_n1031_;
  assign new_n1033_ = ~new_n1032_ & ~new_n1028_ & ~new_n1020_ & ~new_n1024_;
  assign new_n1034_ = ~pi09 & ~new_n22_ & ~pi07;
  assign new_n1035_ = ~new_n1034_ | ~new_n37_ | ~new_n26_ | ~pi14;
  assign new_n1036_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1037_ = ~pi02 | ~pi00;
  assign new_n1038_ = ~new_n1037_ & ~pi03 & ~new_n1035_ & ~new_n1036_;
  assign new_n1039_ = ~new_n22_ & ~pi13 & ~pi09;
  assign new_n1040_ = ~pi14 | ~new_n1039_ | ~new_n37_;
  assign new_n1041_ = ~pi02 | ~new_n66_ | ~new_n24_;
  assign new_n1042_ = ~new_n64_ & ~pi05 & ~new_n1040_ & ~new_n1041_;
  assign new_n1043_ = ~new_n22_ & ~pi13 & ~pi09;
  assign new_n1044_ = ~pi14 | ~new_n1043_ | ~new_n37_;
  assign new_n1045_ = ~pi00 | ~new_n66_ | ~pi02;
  assign new_n1046_ = ~new_n64_ & ~pi05 & ~new_n1044_ & ~new_n1045_;
  assign new_n1047_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1048_ = ~pi04 | ~new_n1047_ | ~pi07;
  assign new_n1049_ = ~pi11 | ~new_n62_ | ~new_n79_;
  assign new_n1050_ = ~new_n26_ & ~pi14 & ~new_n1048_ & ~new_n1049_;
  assign new_n1051_ = ~new_n1050_ & ~new_n1046_ & ~new_n1038_ & ~new_n1042_;
  assign new_n1052_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1053_ = ~pi04 | ~new_n1052_ | ~pi07;
  assign new_n1054_ = ~pi11 | ~new_n26_ | ~new_n79_;
  assign new_n1055_ = ~new_n27_ & ~pi15 & ~new_n1053_ & ~new_n1054_;
  assign new_n1056_ = ~new_n41_ & ~pi03 & ~new_n25_;
  assign new_n1057_ = ~pi04 | ~new_n1056_ | ~pi07;
  assign new_n1058_ = ~pi11 | ~new_n26_ | ~new_n79_;
  assign new_n1059_ = ~new_n27_ & ~pi15 & ~new_n1057_ & ~new_n1058_;
  assign new_n1060_ = ~pi00 & ~new_n24_;
  assign new_n1061_ = ~pi03 | ~new_n1060_ | ~pi07 | ~pi04;
  assign new_n1062_ = ~pi11 | ~new_n62_ | ~new_n79_;
  assign new_n1063_ = ~new_n26_ & ~pi14 & ~new_n1061_ & ~new_n1062_;
  assign new_n1064_ = ~pi09 & ~new_n22_ & ~pi07;
  assign new_n1065_ = ~new_n1064_ | ~new_n27_ | ~new_n62_ | ~pi13;
  assign new_n1066_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1067_ = ~new_n41_ | ~pi01;
  assign new_n1068_ = ~new_n1067_ & ~pi02 & ~new_n1065_ & ~new_n1066_;
  assign new_n1069_ = ~new_n1068_ & ~new_n1063_ & ~new_n1055_ & ~new_n1059_;
  assign new_n1070_ = ~new_n1002_ | ~new_n1033_ | ~new_n1051_ | ~new_n1069_;
  assign new_n1071_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1072_ = ~pi04 | ~new_n1071_ | ~pi07;
  assign new_n1073_ = ~pi11 | ~new_n62_ | ~new_n79_;
  assign new_n1074_ = ~new_n26_ & ~pi14 & ~new_n1072_ & ~new_n1073_;
  assign new_n1075_ = ~new_n41_ & ~pi03 & ~new_n25_;
  assign new_n1076_ = ~pi04 | ~new_n1075_ | ~pi07;
  assign new_n1077_ = ~pi11 | ~new_n62_ | ~new_n79_;
  assign new_n1078_ = ~new_n26_ & ~pi14 & ~new_n1076_ & ~new_n1077_;
  assign new_n1079_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1080_ = ~new_n1079_ | ~new_n89_ | ~pi07 | ~pi04;
  assign new_n1081_ = ~pi12 | ~new_n37_ | ~pi14;
  assign new_n1082_ = ~pi09 | ~pi10;
  assign new_n1083_ = ~new_n1082_ & ~pi11 & ~new_n1080_ & ~new_n1081_;
  assign new_n1084_ = ~new_n24_ & ~new_n66_ & ~pi00;
  assign new_n1085_ = ~new_n1084_ | ~new_n89_ | ~pi07 | ~pi04;
  assign new_n1086_ = ~pi12 | ~new_n37_ | ~pi14;
  assign new_n1087_ = ~pi09 | ~pi10;
  assign new_n1088_ = ~new_n1087_ & ~pi11 & ~new_n1085_ & ~new_n1086_;
  assign new_n1089_ = ~new_n1088_ & ~new_n1083_ & ~new_n1074_ & ~new_n1078_;
  assign new_n1090_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1091_ = ~new_n62_ & ~new_n27_ & ~new_n1090_ & ~pi15;
  assign new_n1092_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1093_ = ~pi06 & ~pi08 & ~pi05;
  assign new_n1094_ = ~new_n1093_ | ~new_n1091_ | ~new_n1092_;
  assign new_n1095_ = ~new_n89_ | ~pi09 | ~new_n22_ | ~pi10;
  assign new_n1096_ = ~new_n62_ & ~new_n27_ & ~new_n1095_ & ~pi15;
  assign new_n1097_ = ~pi04 & ~pi02 & ~pi00 & ~new_n24_;
  assign new_n1098_ = ~new_n104_ & ~pi07 & ~new_n57_;
  assign new_n1099_ = ~new_n1098_ | ~new_n1096_ | ~new_n1097_;
  assign new_n1100_ = ~new_n89_ | ~pi09 | ~new_n22_ | ~pi10;
  assign new_n1101_ = ~new_n62_ & ~new_n27_ & ~new_n1100_ & ~pi15;
  assign new_n1102_ = ~new_n66_ & ~pi04 & ~pi00 & ~new_n24_;
  assign new_n1103_ = ~new_n104_ & ~pi07 & ~new_n57_;
  assign new_n1104_ = ~new_n1103_ | ~new_n1101_ | ~new_n1102_;
  assign new_n1105_ = ~new_n1089_ | ~new_n1094_ | ~new_n1099_ | ~new_n1104_;
  assign new_n1106_ = ~new_n24_ | ~pi02;
  assign new_n1107_ = ~pi06 & ~pi05 & ~pi03 & ~new_n1106_;
  assign new_n1108_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1109_ = ~new_n1107_ | ~new_n1108_ | ~new_n27_ | ~pi13;
  assign new_n1110_ = ~pi02 | ~pi00;
  assign new_n1111_ = ~pi06 & ~pi05 & ~pi03 & ~new_n1110_;
  assign new_n1112_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1113_ = ~new_n1111_ | ~new_n1112_ | ~new_n27_ | ~pi13;
  assign new_n1114_ = ~new_n57_ | ~pi04;
  assign new_n1115_ = ~new_n25_ & ~pi01 & ~new_n1114_ & ~pi03;
  assign new_n1116_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1117_ = ~new_n1115_ | ~new_n1116_ | ~new_n27_ | ~pi13;
  assign new_n1118_ = ~pi02 | ~pi00;
  assign new_n1119_ = ~new_n56_ & ~pi06 & ~pi03 & ~new_n1118_;
  assign new_n1120_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1121_ = ~new_n1119_ | ~new_n1120_ | ~new_n27_ | ~pi13;
  assign new_n1122_ = ~new_n1109_ | ~new_n1113_ | ~new_n1117_ | ~new_n1121_;
  assign new_n1123_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1124_ = ~new_n25_ & ~pi01 & ~new_n1123_ & ~pi03;
  assign new_n1125_ = ~new_n26_ & ~pi14 & ~pi12;
  assign new_n1126_ = ~pi07 & ~pi09;
  assign new_n1127_ = ~new_n1124_ | ~new_n1125_ | ~pi11 | ~new_n1126_;
  assign new_n1128_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1129_ = ~new_n41_ & ~new_n25_ & ~new_n1128_ & ~pi03;
  assign new_n1130_ = ~new_n26_ & ~pi14 & ~pi12;
  assign new_n1131_ = ~pi07 & ~pi09;
  assign new_n1132_ = ~new_n1129_ | ~new_n1130_ | ~pi11 | ~new_n1131_;
  assign new_n1133_ = ~new_n104_ | ~pi07;
  assign new_n1134_ = ~new_n25_ & ~pi01 & ~new_n1133_ & ~pi03;
  assign new_n1135_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1136_ = ~new_n1134_ | ~new_n1135_ | ~new_n27_ | ~pi13;
  assign new_n1137_ = ~pi02 | ~pi00;
  assign new_n1138_ = ~new_n64_ & ~pi05 & ~pi03 & ~new_n1137_;
  assign new_n1139_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1140_ = ~new_n1138_ | ~new_n1139_ | ~new_n27_ | ~pi13;
  assign new_n1141_ = ~new_n1127_ | ~new_n1132_ | ~new_n1136_ | ~new_n1140_;
  assign new_n1142_ = ~new_n1141_ & ~new_n1105_ & ~new_n1122_;
  assign new_n1143_ = ~pi00 | ~new_n66_ | ~pi02;
  assign new_n1144_ = ~new_n56_ & ~pi06 & ~new_n1143_ & ~pi08;
  assign new_n1145_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1146_ = ~new_n62_ & ~new_n27_ & ~new_n1145_ & ~pi15;
  assign new_n1147_ = ~new_n1144_ | ~new_n1146_;
  assign new_n1148_ = ~new_n89_ | ~pi09 | ~new_n22_ | ~pi10;
  assign new_n1149_ = ~new_n62_ & ~new_n27_ & ~new_n1148_ & ~pi15;
  assign new_n1150_ = ~pi04 & ~pi03 & ~pi01 & ~new_n25_;
  assign new_n1151_ = ~new_n104_ & ~pi07 & ~new_n57_;
  assign new_n1152_ = ~new_n1151_ | ~new_n1149_ | ~new_n1150_;
  assign new_n1153_ = ~new_n89_ | ~pi09 | ~new_n22_ | ~pi10;
  assign new_n1154_ = ~new_n62_ & ~new_n27_ & ~new_n1153_ & ~pi15;
  assign new_n1155_ = ~pi04 & ~pi03 & ~new_n25_ & ~new_n41_;
  assign new_n1156_ = ~new_n104_ & ~pi07 & ~new_n57_;
  assign new_n1157_ = ~new_n1156_ | ~new_n1154_ | ~new_n1155_;
  assign new_n1158_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1159_ = ~new_n62_ & ~new_n27_ & ~new_n1158_ & ~pi15;
  assign new_n1160_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1161_ = ~new_n64_ & ~pi08 & ~pi05;
  assign new_n1162_ = ~new_n1161_ | ~new_n1159_ | ~new_n1160_;
  assign new_n1163_ = ~new_n1147_ | ~new_n1152_ | ~new_n1157_ | ~new_n1162_;
  assign new_n1164_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1165_ = ~new_n1164_ | ~new_n89_ | ~pi07 | ~pi04;
  assign new_n1166_ = ~pi12 | ~new_n37_ | ~pi14;
  assign new_n1167_ = ~pi09 | ~pi10;
  assign new_n1168_ = ~new_n1167_ & ~pi11 & ~new_n1165_ & ~new_n1166_;
  assign new_n1169_ = ~new_n64_ & ~pi08 & ~pi05;
  assign new_n1170_ = ~new_n1169_ | ~new_n66_ | ~pi02 | ~pi00;
  assign new_n1171_ = ~pi12 | ~new_n37_ | ~pi14;
  assign new_n1172_ = ~pi09 | ~pi10;
  assign new_n1173_ = ~new_n1172_ & ~pi11 & ~new_n1170_ & ~new_n1171_;
  assign new_n1174_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1175_ = ~new_n1174_ | ~new_n89_ | ~pi07 | ~pi04;
  assign new_n1176_ = ~pi14 | ~new_n37_ | ~new_n26_;
  assign new_n1177_ = ~pi09 | ~pi10;
  assign new_n1178_ = ~new_n1177_ & ~pi11 & ~new_n1175_ & ~new_n1176_;
  assign new_n1179_ = ~new_n1178_ & ~new_n1173_ & ~new_n1163_ & ~new_n1168_;
  assign new_n1180_ = ~pi06 & ~pi08 & ~pi05;
  assign new_n1181_ = ~new_n1180_ | ~pi03 | ~new_n41_ | ~pi01;
  assign new_n1182_ = ~pi12 | ~new_n37_ | ~pi14;
  assign new_n1183_ = ~pi09 | ~pi10;
  assign new_n1184_ = ~new_n1183_ & ~pi11 & ~new_n1181_ & ~new_n1182_;
  assign new_n1185_ = ~new_n56_ & ~pi08 & ~pi06;
  assign new_n1186_ = ~new_n1185_ | ~new_n25_ | ~new_n41_ | ~pi01;
  assign new_n1187_ = ~pi12 | ~new_n37_ | ~pi14;
  assign new_n1188_ = ~pi09 | ~pi10;
  assign new_n1189_ = ~new_n1188_ & ~pi11 & ~new_n1186_ & ~new_n1187_;
  assign new_n1190_ = ~new_n56_ & ~pi08 & ~pi06;
  assign new_n1191_ = ~new_n1190_ | ~pi03 | ~new_n41_ | ~pi01;
  assign new_n1192_ = ~pi12 | ~new_n37_ | ~pi14;
  assign new_n1193_ = ~pi09 | ~pi10;
  assign new_n1194_ = ~new_n1193_ & ~pi11 & ~new_n1191_ & ~new_n1192_;
  assign new_n1195_ = ~new_n64_ & ~pi08 & ~pi05;
  assign new_n1196_ = ~new_n1195_ | ~new_n25_ | ~new_n41_ | ~pi01;
  assign new_n1197_ = ~pi12 | ~new_n37_ | ~pi14;
  assign new_n1198_ = ~pi09 | ~pi10;
  assign new_n1199_ = ~new_n1198_ & ~pi11 & ~new_n1196_ & ~new_n1197_;
  assign new_n1200_ = ~new_n1199_ & ~new_n1194_ & ~new_n1184_ & ~new_n1189_;
  assign new_n1201_ = ~new_n64_ & ~pi08 & ~pi05;
  assign new_n1202_ = ~new_n1201_ | ~pi03 | ~new_n41_ | ~pi01;
  assign new_n1203_ = ~pi12 | ~new_n37_ | ~pi14;
  assign new_n1204_ = ~pi09 | ~pi10;
  assign new_n1205_ = ~new_n1204_ & ~pi11 & ~new_n1202_ & ~new_n1203_;
  assign new_n1206_ = ~pi06 & ~pi08 & ~pi05;
  assign new_n1207_ = ~new_n1206_ | ~new_n66_ | ~new_n24_ | ~pi02;
  assign new_n1208_ = ~pi12 | ~new_n37_ | ~pi14;
  assign new_n1209_ = ~pi09 | ~pi10;
  assign new_n1210_ = ~new_n1209_ & ~pi11 & ~new_n1207_ & ~new_n1208_;
  assign new_n1211_ = ~pi06 & ~pi08 & ~pi05;
  assign new_n1212_ = ~new_n1211_ | ~new_n66_ | ~pi02 | ~pi00;
  assign new_n1213_ = ~pi12 | ~new_n37_ | ~pi14;
  assign new_n1214_ = ~pi09 | ~pi10;
  assign new_n1215_ = ~new_n1214_ & ~pi11 & ~new_n1212_ & ~new_n1213_;
  assign new_n1216_ = ~new_n56_ & ~pi08 & ~pi06;
  assign new_n1217_ = ~new_n1216_ | ~new_n66_ | ~new_n24_ | ~pi02;
  assign new_n1218_ = ~pi12 | ~new_n37_ | ~pi14;
  assign new_n1219_ = ~pi09 | ~pi10;
  assign new_n1220_ = ~new_n1219_ & ~pi11 & ~new_n1217_ & ~new_n1218_;
  assign new_n1221_ = ~new_n1220_ & ~new_n1215_ & ~new_n1205_ & ~new_n1210_;
  assign new_n1222_ = ~new_n1142_ | ~new_n1179_ | ~new_n1200_ | ~new_n1221_;
  assign new_n1223_ = ~new_n89_ | ~pi09 | ~new_n22_ | ~pi10;
  assign new_n1224_ = ~new_n27_ & ~pi13 & ~new_n1223_ & ~pi15;
  assign new_n1225_ = ~pi04 & ~pi03 & ~new_n25_ & ~new_n41_;
  assign new_n1226_ = ~new_n104_ & ~pi07 & ~new_n57_;
  assign new_n1227_ = ~new_n1226_ | ~new_n1224_ | ~new_n1225_;
  assign new_n1228_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1229_ = ~new_n27_ & ~pi13 & ~new_n1228_ & ~pi15;
  assign new_n1230_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1231_ = ~new_n64_ & ~pi08 & ~pi05;
  assign new_n1232_ = ~new_n1231_ | ~new_n1229_ | ~new_n1230_;
  assign new_n1233_ = ~pi00 | ~new_n66_ | ~pi02;
  assign new_n1234_ = ~new_n64_ & ~pi05 & ~new_n1233_ & ~pi08;
  assign new_n1235_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1236_ = ~new_n27_ & ~pi13 & ~new_n1235_ & ~pi15;
  assign new_n1237_ = ~new_n1234_ | ~new_n1236_;
  assign new_n1238_ = ~pi04 | ~new_n89_ | ~pi07;
  assign new_n1239_ = ~new_n25_ & ~pi01 & ~new_n1238_ & ~pi03;
  assign new_n1240_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1241_ = ~new_n27_ & ~pi13 & ~new_n1240_ & ~pi15;
  assign new_n1242_ = ~new_n1239_ | ~new_n1241_;
  assign new_n1243_ = ~new_n1227_ | ~new_n1232_ | ~new_n1237_ | ~new_n1242_;
  assign new_n1244_ = ~pi04 | ~new_n89_ | ~pi07;
  assign new_n1245_ = ~new_n41_ & ~new_n25_ & ~new_n1244_ & ~pi03;
  assign new_n1246_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1247_ = ~new_n27_ & ~pi13 & ~new_n1246_ & ~pi15;
  assign new_n1248_ = ~new_n1245_ | ~new_n1247_;
  assign new_n1249_ = ~pi08 | ~pi11;
  assign new_n1250_ = ~new_n37_ & ~new_n26_ & ~pi12 & ~new_n1249_;
  assign new_n1251_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1252_ = ~new_n1250_ | ~new_n1251_ | ~pi07 | ~pi04;
  assign new_n1253_ = ~pi08 | ~pi11;
  assign new_n1254_ = ~new_n37_ & ~new_n26_ & ~pi12 & ~new_n1253_;
  assign new_n1255_ = ~new_n24_ & ~new_n66_ & ~pi00;
  assign new_n1256_ = ~new_n1254_ | ~new_n1255_ | ~pi07 | ~pi04;
  assign new_n1257_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1258_ = ~new_n24_ & ~pi00 & ~new_n1257_ & ~pi02;
  assign new_n1259_ = ~pi08 | ~pi11 | ~new_n64_;
  assign new_n1260_ = ~new_n26_ & ~pi12 & ~new_n1259_ & ~new_n37_;
  assign new_n1261_ = ~new_n1258_ | ~new_n1260_;
  assign new_n1262_ = ~new_n1248_ | ~new_n1252_ | ~new_n1256_ | ~new_n1261_;
  assign new_n1263_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1264_ = ~new_n24_ & ~pi00 & ~new_n1263_ & ~new_n66_;
  assign new_n1265_ = ~pi08 | ~pi11 | ~new_n64_;
  assign new_n1266_ = ~new_n26_ & ~pi12 & ~new_n1265_ & ~new_n37_;
  assign new_n1267_ = ~new_n1264_ | ~new_n1266_;
  assign new_n1268_ = ~new_n41_ | ~pi01;
  assign new_n1269_ = ~pi06 & ~pi05 & ~pi02 & ~new_n1268_;
  assign new_n1270_ = ~new_n22_ & ~pi12 & ~new_n89_;
  assign new_n1271_ = ~new_n1269_ | ~new_n1270_ | ~pi13 | ~pi15;
  assign new_n1272_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1273_ = ~pi06 & ~new_n1272_ & ~pi05;
  assign new_n1274_ = ~new_n22_ & ~pi12 & ~new_n89_;
  assign new_n1275_ = ~new_n1273_ | ~new_n1274_ | ~pi13 | ~pi15;
  assign new_n1276_ = ~pi08 | ~pi11;
  assign new_n1277_ = ~new_n37_ & ~new_n26_ & ~pi12 & ~new_n1276_;
  assign new_n1278_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1279_ = ~new_n1277_ | ~new_n1278_ | ~new_n57_ | ~pi04;
  assign new_n1280_ = ~new_n1267_ | ~new_n1271_ | ~new_n1275_ | ~new_n1279_;
  assign new_n1281_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1282_ = ~new_n64_ & ~new_n1281_ & ~pi05;
  assign new_n1283_ = ~new_n22_ & ~pi12 & ~new_n89_;
  assign new_n1284_ = ~new_n1282_ | ~new_n1283_ | ~pi13 | ~pi15;
  assign new_n1285_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1286_ = ~new_n56_ & ~new_n1285_ & ~pi06;
  assign new_n1287_ = ~new_n22_ & ~pi12 & ~new_n89_;
  assign new_n1288_ = ~new_n1286_ | ~new_n1287_ | ~pi13 | ~pi15;
  assign new_n1289_ = ~pi08 | ~pi11;
  assign new_n1290_ = ~new_n37_ & ~new_n26_ & ~pi12 & ~new_n1289_;
  assign new_n1291_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1292_ = ~new_n1290_ | ~new_n1291_ | ~new_n104_ | ~pi07;
  assign new_n1293_ = ~new_n1292_ | ~new_n1284_ | ~new_n1288_;
  assign new_n1294_ = ~new_n1293_ & ~new_n1280_ & ~new_n1243_ & ~new_n1262_;
  assign new_n1295_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1296_ = ~new_n27_ & ~pi13 & ~new_n1295_ & ~pi15;
  assign new_n1297_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1298_ = ~new_n64_ & ~pi08 & ~pi05;
  assign new_n1299_ = ~new_n1298_ | ~new_n1296_ | ~new_n1297_;
  assign new_n1300_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1301_ = ~new_n27_ & ~pi13 & ~new_n1300_ & ~pi15;
  assign new_n1302_ = ~new_n64_ & ~pi08 & ~pi05;
  assign new_n1303_ = ~pi00 & ~new_n24_;
  assign new_n1304_ = ~new_n1301_ | ~new_n1302_ | ~pi03 | ~new_n1303_;
  assign new_n1305_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1306_ = ~new_n27_ & ~pi13 & ~new_n1305_ & ~pi15;
  assign new_n1307_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1308_ = ~pi06 & ~pi08 & ~pi05;
  assign new_n1309_ = ~new_n1308_ | ~new_n1306_ | ~new_n1307_;
  assign new_n1310_ = ~pi00 | ~new_n66_ | ~pi02;
  assign new_n1311_ = ~pi06 & ~pi05 & ~new_n1310_ & ~pi08;
  assign new_n1312_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1313_ = ~new_n27_ & ~pi13 & ~new_n1312_ & ~pi15;
  assign new_n1314_ = ~new_n1311_ | ~new_n1313_;
  assign new_n1315_ = ~new_n1299_ | ~new_n1304_ | ~new_n1309_ | ~new_n1314_;
  assign new_n1316_ = ~pi04 & ~pi03 & ~pi01 & ~new_n25_;
  assign new_n1317_ = ~new_n1316_ | ~new_n64_ | ~pi06 | ~pi05;
  assign new_n1318_ = ~new_n89_ | ~pi09 | ~new_n22_ | ~pi10;
  assign new_n1319_ = ~new_n26_ | ~pi14;
  assign new_n1320_ = ~new_n1319_ & ~pi15 & ~new_n1317_ & ~new_n1318_;
  assign new_n1321_ = ~new_n56_ & ~pi08 & ~pi06;
  assign new_n1322_ = ~new_n1321_ | ~new_n66_ | ~new_n24_ | ~pi02;
  assign new_n1323_ = ~pi14 | ~new_n37_ | ~new_n26_;
  assign new_n1324_ = ~pi09 | ~pi10;
  assign new_n1325_ = ~new_n1324_ & ~pi11 & ~new_n1322_ & ~new_n1323_;
  assign new_n1326_ = ~new_n56_ & ~pi08 & ~pi06;
  assign new_n1327_ = ~new_n1326_ | ~new_n66_ | ~pi02 | ~pi00;
  assign new_n1328_ = ~pi14 | ~new_n37_ | ~new_n26_;
  assign new_n1329_ = ~pi09 | ~pi10;
  assign new_n1330_ = ~new_n1329_ & ~pi11 & ~new_n1327_ & ~new_n1328_;
  assign new_n1331_ = ~new_n1330_ & ~new_n1325_ & ~new_n1315_ & ~new_n1320_;
  assign new_n1332_ = ~new_n41_ & ~pi03 & ~new_n25_;
  assign new_n1333_ = ~new_n1332_ | ~new_n89_ | ~pi07 | ~pi04;
  assign new_n1334_ = ~pi12 | ~new_n37_ | ~pi14;
  assign new_n1335_ = ~pi09 | ~pi10;
  assign new_n1336_ = ~new_n1335_ & ~pi11 & ~new_n1333_ & ~new_n1334_;
  assign new_n1337_ = ~new_n27_ & ~pi15 & ~pi13;
  assign new_n1338_ = ~new_n1337_ | ~new_n22_ | ~pi09 | ~pi10;
  assign new_n1339_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1340_ = ~pi07 | ~pi04;
  assign new_n1341_ = ~new_n1340_ & ~pi08 & ~new_n1338_ & ~new_n1339_;
  assign new_n1342_ = ~pi04 & ~pi02 & ~pi00 & ~new_n24_;
  assign new_n1343_ = ~new_n1342_ | ~new_n64_ | ~pi06 | ~pi05;
  assign new_n1344_ = ~new_n89_ | ~pi09 | ~new_n22_ | ~pi10;
  assign new_n1345_ = ~new_n26_ | ~pi14;
  assign new_n1346_ = ~new_n1345_ & ~pi15 & ~new_n1343_ & ~new_n1344_;
  assign new_n1347_ = ~new_n19_ & ~pi11 & ~pi08 & ~new_n79_;
  assign new_n1348_ = ~new_n1347_ | ~new_n37_ | ~new_n26_ | ~pi14;
  assign new_n1349_ = ~new_n41_ | ~pi01 | ~new_n56_ | ~pi03;
  assign new_n1350_ = ~pi06 | ~pi05;
  assign new_n1351_ = ~new_n1350_ & ~pi07 & ~new_n1348_ & ~new_n1349_;
  assign new_n1352_ = ~new_n1351_ & ~new_n1346_ & ~new_n1336_ & ~new_n1341_;
  assign new_n1353_ = ~pi06 & ~pi08 & ~pi05;
  assign new_n1354_ = ~new_n1353_ | ~new_n25_ | ~new_n41_ | ~pi01;
  assign new_n1355_ = ~pi14 | ~new_n37_ | ~new_n26_;
  assign new_n1356_ = ~pi09 | ~pi10;
  assign new_n1357_ = ~new_n1356_ & ~pi11 & ~new_n1354_ & ~new_n1355_;
  assign new_n1358_ = ~pi06 & ~pi08 & ~pi05;
  assign new_n1359_ = ~new_n1358_ | ~pi03 | ~new_n41_ | ~pi01;
  assign new_n1360_ = ~pi14 | ~new_n37_ | ~new_n26_;
  assign new_n1361_ = ~pi09 | ~pi10;
  assign new_n1362_ = ~new_n1361_ & ~pi11 & ~new_n1359_ & ~new_n1360_;
  assign new_n1363_ = ~new_n56_ & ~pi08 & ~pi06;
  assign new_n1364_ = ~new_n1363_ | ~new_n25_ | ~new_n41_ | ~pi01;
  assign new_n1365_ = ~pi14 | ~new_n37_ | ~new_n26_;
  assign new_n1366_ = ~pi09 | ~pi10;
  assign new_n1367_ = ~new_n1366_ & ~pi11 & ~new_n1364_ & ~new_n1365_;
  assign new_n1368_ = ~new_n56_ & ~pi08 & ~pi06;
  assign new_n1369_ = ~new_n1368_ | ~pi03 | ~new_n41_ | ~pi01;
  assign new_n1370_ = ~pi14 | ~new_n37_ | ~new_n26_;
  assign new_n1371_ = ~pi09 | ~pi10;
  assign new_n1372_ = ~new_n1371_ & ~pi11 & ~new_n1369_ & ~new_n1370_;
  assign new_n1373_ = ~new_n1372_ & ~new_n1367_ & ~new_n1357_ & ~new_n1362_;
  assign new_n1374_ = ~new_n1294_ | ~new_n1331_ | ~new_n1352_ | ~new_n1373_;
  assign new_n1375_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1376_ = ~pi06 & ~new_n1375_ & ~pi05;
  assign new_n1377_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1378_ = ~new_n1376_ | ~new_n1377_ | ~pi13 | ~pi15;
  assign new_n1379_ = ~pi13 | ~pi15;
  assign new_n1380_ = ~new_n89_ & ~pi10 & ~new_n1379_ & ~pi12;
  assign new_n1381_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1382_ = ~new_n1380_ | ~new_n1381_ | ~new_n57_ | ~pi04;
  assign new_n1383_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1384_ = ~new_n56_ & ~new_n1383_ & ~pi06;
  assign new_n1385_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1386_ = ~new_n1384_ | ~new_n1385_ | ~pi13 | ~pi15;
  assign new_n1387_ = ~pi13 | ~pi15;
  assign new_n1388_ = ~new_n89_ & ~pi10 & ~new_n1387_ & ~pi12;
  assign new_n1389_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1390_ = ~new_n1388_ | ~new_n1389_ | ~new_n104_ | ~pi07;
  assign new_n1391_ = ~new_n1378_ | ~new_n1382_ | ~new_n1386_ | ~new_n1390_;
  assign new_n1392_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1393_ = ~new_n64_ & ~new_n1392_ & ~pi05;
  assign new_n1394_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1395_ = ~new_n1393_ | ~new_n1394_ | ~pi13 | ~pi15;
  assign new_n1396_ = ~new_n24_ | ~pi02;
  assign new_n1397_ = ~pi06 & ~pi05 & ~pi03 & ~new_n1396_;
  assign new_n1398_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1399_ = ~new_n1397_ | ~new_n1398_ | ~pi13 | ~pi15;
  assign new_n1400_ = ~pi02 | ~pi00;
  assign new_n1401_ = ~pi06 & ~pi05 & ~pi03 & ~new_n1400_;
  assign new_n1402_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1403_ = ~new_n1401_ | ~new_n1402_ | ~pi13 | ~pi15;
  assign new_n1404_ = ~pi13 | ~pi15;
  assign new_n1405_ = ~new_n89_ & ~pi10 & ~new_n1404_ & ~pi12;
  assign new_n1406_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1407_ = ~new_n1405_ | ~new_n1406_ | ~new_n57_ | ~pi04;
  assign new_n1408_ = ~new_n1395_ | ~new_n1399_ | ~new_n1403_ | ~new_n1407_;
  assign new_n1409_ = ~pi02 | ~pi00;
  assign new_n1410_ = ~new_n56_ & ~pi06 & ~pi03 & ~new_n1409_;
  assign new_n1411_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1412_ = ~new_n1410_ | ~new_n1411_ | ~pi13 | ~pi15;
  assign new_n1413_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1414_ = ~new_n25_ & ~pi01 & ~new_n1413_ & ~pi03;
  assign new_n1415_ = ~new_n89_ & ~pi10 & ~pi07;
  assign new_n1416_ = ~pi12 & ~new_n26_;
  assign new_n1417_ = ~new_n1414_ | ~new_n1415_ | ~pi15 | ~new_n1416_;
  assign new_n1418_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1419_ = ~new_n41_ & ~new_n25_ & ~new_n1418_ & ~pi03;
  assign new_n1420_ = ~new_n89_ & ~pi10 & ~pi07;
  assign new_n1421_ = ~pi12 & ~new_n26_;
  assign new_n1422_ = ~new_n1419_ | ~new_n1420_ | ~pi15 | ~new_n1421_;
  assign new_n1423_ = ~pi13 | ~pi15;
  assign new_n1424_ = ~new_n89_ & ~pi10 & ~new_n1423_ & ~pi12;
  assign new_n1425_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1426_ = ~new_n1424_ | ~new_n1425_ | ~new_n104_ | ~pi07;
  assign new_n1427_ = ~new_n1412_ | ~new_n1417_ | ~new_n1422_ | ~new_n1426_;
  assign new_n1428_ = ~pi13 | ~pi15;
  assign new_n1429_ = ~new_n89_ & ~pi10 & ~new_n1428_ & ~pi12;
  assign new_n1430_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1431_ = ~new_n1429_ | ~new_n1430_ | ~pi07 | ~pi04;
  assign new_n1432_ = ~pi02 | ~pi00;
  assign new_n1433_ = ~new_n64_ & ~pi05 & ~pi03 & ~new_n1432_;
  assign new_n1434_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1435_ = ~new_n1433_ | ~new_n1434_ | ~pi13 | ~pi15;
  assign new_n1436_ = ~pi13 | ~pi15;
  assign new_n1437_ = ~pi10 & ~pi09 & ~new_n1436_ & ~pi12;
  assign new_n1438_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1439_ = ~new_n1437_ | ~new_n1438_ | ~pi07 | ~pi04;
  assign new_n1440_ = ~new_n1439_ | ~new_n1431_ | ~new_n1435_;
  assign new_n1441_ = ~new_n1440_ & ~new_n1427_ & ~new_n1391_ & ~new_n1408_;
  assign new_n1442_ = ~pi13 | ~pi15;
  assign new_n1443_ = ~new_n89_ & ~pi10 & ~new_n1442_ & ~pi12;
  assign new_n1444_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1445_ = ~new_n1443_ | ~new_n1444_ | ~pi07 | ~pi04;
  assign new_n1446_ = ~pi08 | ~pi11;
  assign new_n1447_ = ~new_n37_ & ~new_n26_ & ~pi12 & ~new_n1446_;
  assign new_n1448_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1449_ = ~new_n1447_ | ~new_n1448_ | ~pi07 | ~pi04;
  assign new_n1450_ = ~pi08 | ~pi11;
  assign new_n1451_ = ~new_n37_ & ~new_n26_ & ~pi12 & ~new_n1450_;
  assign new_n1452_ = ~new_n41_ & ~pi03 & ~new_n25_;
  assign new_n1453_ = ~new_n1451_ | ~new_n1452_ | ~pi07 | ~pi04;
  assign new_n1454_ = ~pi13 | ~pi15;
  assign new_n1455_ = ~new_n89_ & ~pi10 & ~new_n1454_ & ~pi12;
  assign new_n1456_ = ~new_n24_ & ~new_n66_ & ~pi00;
  assign new_n1457_ = ~new_n1455_ | ~new_n1456_ | ~pi07 | ~pi04;
  assign new_n1458_ = ~new_n1445_ | ~new_n1449_ | ~new_n1453_ | ~new_n1457_;
  assign new_n1459_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1460_ = ~pi15 | ~new_n1459_ | ~pi13;
  assign new_n1461_ = ~pi01 | ~new_n25_ | ~new_n41_;
  assign new_n1462_ = ~pi06 & ~pi05 & ~new_n1460_ & ~new_n1461_;
  assign new_n1463_ = ~new_n89_ & ~pi10 & ~pi07;
  assign new_n1464_ = ~new_n1463_ | ~pi15 | ~new_n62_ | ~pi13;
  assign new_n1465_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1466_ = ~new_n41_ | ~pi01;
  assign new_n1467_ = ~new_n1466_ & ~pi02 & ~new_n1464_ & ~new_n1465_;
  assign new_n1468_ = ~new_n89_ & ~pi10 & ~pi07;
  assign new_n1469_ = ~new_n1468_ | ~pi15 | ~new_n62_ | ~pi13;
  assign new_n1470_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1471_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1472_ = ~new_n1471_ & ~new_n1469_ & ~new_n1470_;
  assign new_n1473_ = ~new_n1472_ & ~new_n1467_ & ~new_n1458_ & ~new_n1462_;
  assign new_n1474_ = ~new_n22_ & ~pi12 & ~new_n89_;
  assign new_n1475_ = ~pi15 | ~new_n1474_ | ~pi13;
  assign new_n1476_ = ~pi02 | ~new_n66_ | ~new_n24_;
  assign new_n1477_ = ~pi06 & ~pi05 & ~new_n1475_ & ~new_n1476_;
  assign new_n1478_ = ~new_n22_ & ~pi12 & ~new_n89_;
  assign new_n1479_ = ~pi15 | ~new_n1478_ | ~pi13;
  assign new_n1480_ = ~pi00 | ~new_n66_ | ~pi02;
  assign new_n1481_ = ~pi06 & ~pi05 & ~new_n1479_ & ~new_n1480_;
  assign new_n1482_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1483_ = ~pi04 | ~new_n1482_ | ~new_n57_;
  assign new_n1484_ = ~pi11 | ~new_n62_ | ~pi08;
  assign new_n1485_ = ~new_n37_ & ~new_n26_ & ~new_n1483_ & ~new_n1484_;
  assign new_n1486_ = ~new_n22_ & ~pi12 & ~new_n89_;
  assign new_n1487_ = ~pi15 | ~new_n1486_ | ~pi13;
  assign new_n1488_ = ~pi00 | ~new_n66_ | ~pi02;
  assign new_n1489_ = ~new_n56_ & ~pi06 & ~new_n1487_ & ~new_n1488_;
  assign new_n1490_ = ~new_n1489_ & ~new_n1485_ & ~new_n1477_ & ~new_n1481_;
  assign new_n1491_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1492_ = ~new_n1491_ | ~pi06 | ~new_n56_ | ~pi05;
  assign new_n1493_ = ~pi08 | ~pi11 | ~new_n64_;
  assign new_n1494_ = ~pi13 | ~pi15 | ~new_n62_;
  assign new_n1495_ = ~new_n1494_ & ~new_n1492_ & ~new_n1493_;
  assign new_n1496_ = ~pi00 | ~new_n66_ | ~pi02;
  assign new_n1497_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1498_ = ~pi08 | ~pi11 | ~new_n64_;
  assign new_n1499_ = ~pi13 | ~pi15 | ~new_n62_;
  assign new_n1500_ = ~new_n1499_ & ~new_n1498_ & ~new_n1496_ & ~new_n1497_;
  assign new_n1501_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1502_ = ~pi07 | ~new_n1501_ | ~new_n104_;
  assign new_n1503_ = ~pi11 | ~new_n62_ | ~pi08;
  assign new_n1504_ = ~new_n37_ & ~new_n26_ & ~new_n1502_ & ~new_n1503_;
  assign new_n1505_ = ~new_n22_ & ~pi12 & ~new_n89_;
  assign new_n1506_ = ~pi15 | ~new_n1505_ | ~pi13;
  assign new_n1507_ = ~pi00 | ~new_n66_ | ~pi02;
  assign new_n1508_ = ~new_n64_ & ~pi05 & ~new_n1506_ & ~new_n1507_;
  assign new_n1509_ = ~new_n1508_ & ~new_n1504_ & ~new_n1495_ & ~new_n1500_;
  assign new_n1510_ = ~new_n1441_ | ~new_n1473_ | ~new_n1490_ | ~new_n1509_;
  assign new_n1511_ = ~new_n1510_ & ~new_n1374_ & ~new_n1070_ & ~new_n1222_;
  assign new_n1512_ = ~pi13 | ~pi15 | ~new_n62_;
  assign new_n1513_ = ~pi09 & ~pi07 & ~new_n1512_ & ~pi10;
  assign new_n1514_ = ~new_n41_ & ~pi03 & ~new_n25_;
  assign new_n1515_ = ~pi04 & ~new_n104_;
  assign new_n1516_ = ~new_n1513_ | ~new_n1514_ | ~pi06 | ~new_n1515_;
  assign new_n1517_ = ~pi13 | ~pi15;
  assign new_n1518_ = ~pi10 & ~pi09 & ~new_n1517_ & ~pi12;
  assign new_n1519_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1520_ = ~new_n1518_ | ~new_n1519_ | ~new_n104_ | ~pi07;
  assign new_n1521_ = ~pi02 | ~pi00;
  assign new_n1522_ = ~new_n64_ & ~pi05 & ~pi03 & ~new_n1521_;
  assign new_n1523_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n1524_ = ~new_n1522_ | ~new_n1523_ | ~pi13 | ~pi15;
  assign new_n1525_ = ~pi13 | ~pi15;
  assign new_n1526_ = ~pi10 & ~pi09 & ~new_n1525_ & ~pi12;
  assign new_n1527_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1528_ = ~new_n1526_ | ~new_n1527_ | ~pi07 | ~pi04;
  assign new_n1529_ = ~new_n1516_ | ~new_n1520_ | ~new_n1524_ | ~new_n1528_;
  assign new_n1530_ = ~pi13 | ~pi15;
  assign new_n1531_ = ~pi10 & ~pi09 & ~new_n1530_ & ~pi12;
  assign new_n1532_ = ~new_n41_ & ~pi03 & ~new_n25_;
  assign new_n1533_ = ~new_n1531_ | ~new_n1532_ | ~pi07 | ~pi04;
  assign new_n1534_ = ~pi13 | ~pi15;
  assign new_n1535_ = ~new_n22_ & ~pi09 & ~new_n1534_ & ~pi12;
  assign new_n1536_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1537_ = ~new_n1535_ | ~new_n1536_ | ~pi07 | ~pi04;
  assign new_n1538_ = ~pi13 | ~pi15;
  assign new_n1539_ = ~new_n22_ & ~pi09 & ~new_n1538_ & ~pi12;
  assign new_n1540_ = ~new_n24_ & ~new_n66_ & ~pi00;
  assign new_n1541_ = ~new_n1539_ | ~new_n1540_ | ~pi07 | ~pi04;
  assign new_n1542_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1543_ = ~new_n24_ & ~pi00 & ~new_n1542_ & ~pi02;
  assign new_n1544_ = ~new_n26_ & ~new_n37_ & ~pi12;
  assign new_n1545_ = ~pi07 & ~pi09;
  assign new_n1546_ = ~new_n1543_ | ~new_n1544_ | ~pi11 | ~new_n1545_;
  assign new_n1547_ = ~new_n1533_ | ~new_n1537_ | ~new_n1541_ | ~new_n1546_;
  assign new_n1548_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1549_ = ~new_n24_ & ~pi00 & ~new_n1548_ & ~new_n66_;
  assign new_n1550_ = ~new_n26_ & ~new_n37_ & ~pi12;
  assign new_n1551_ = ~pi07 & ~pi09;
  assign new_n1552_ = ~new_n1549_ | ~new_n1550_ | ~pi11 | ~new_n1551_;
  assign new_n1553_ = ~new_n41_ | ~pi01;
  assign new_n1554_ = ~pi06 & ~pi05 & ~pi02 & ~new_n1553_;
  assign new_n1555_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1556_ = ~new_n1554_ | ~new_n1555_ | ~pi13 | ~pi15;
  assign new_n1557_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1558_ = ~pi06 & ~new_n1557_ & ~pi05;
  assign new_n1559_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1560_ = ~new_n1558_ | ~new_n1559_ | ~pi13 | ~pi15;
  assign new_n1561_ = ~pi13 | ~pi15;
  assign new_n1562_ = ~new_n22_ & ~pi09 & ~new_n1561_ & ~pi12;
  assign new_n1563_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1564_ = ~new_n1562_ | ~new_n1563_ | ~new_n57_ | ~pi04;
  assign new_n1565_ = ~new_n1552_ | ~new_n1556_ | ~new_n1560_ | ~new_n1564_;
  assign new_n1566_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1567_ = ~new_n64_ & ~new_n1566_ & ~pi05;
  assign new_n1568_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1569_ = ~new_n1567_ | ~new_n1568_ | ~pi13 | ~pi15;
  assign new_n1570_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1571_ = ~new_n56_ & ~new_n1570_ & ~pi06;
  assign new_n1572_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1573_ = ~new_n1571_ | ~new_n1572_ | ~pi13 | ~pi15;
  assign new_n1574_ = ~pi13 | ~pi15;
  assign new_n1575_ = ~new_n22_ & ~pi09 & ~new_n1574_ & ~pi12;
  assign new_n1576_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1577_ = ~new_n1575_ | ~new_n1576_ | ~new_n104_ | ~pi07;
  assign new_n1578_ = ~new_n1577_ | ~new_n1569_ | ~new_n1573_;
  assign new_n1579_ = ~new_n1578_ & ~new_n1565_ & ~new_n1529_ & ~new_n1547_;
  assign new_n1580_ = ~pi13 | ~pi15;
  assign new_n1581_ = ~pi10 & ~pi09 & ~new_n1580_ & ~pi12;
  assign new_n1582_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1583_ = ~new_n1581_ | ~new_n1582_ | ~new_n104_ | ~pi07;
  assign new_n1584_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1585_ = ~new_n64_ & ~new_n1584_ & ~pi05;
  assign new_n1586_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n1587_ = ~new_n1585_ | ~new_n1586_ | ~pi13 | ~pi15;
  assign new_n1588_ = ~new_n24_ | ~pi02;
  assign new_n1589_ = ~pi06 & ~pi05 & ~pi03 & ~new_n1588_;
  assign new_n1590_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n1591_ = ~new_n1589_ | ~new_n1590_ | ~pi13 | ~pi15;
  assign new_n1592_ = ~pi02 | ~pi00;
  assign new_n1593_ = ~pi06 & ~pi05 & ~pi03 & ~new_n1592_;
  assign new_n1594_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n1595_ = ~new_n1593_ | ~new_n1594_ | ~pi13 | ~pi15;
  assign new_n1596_ = ~new_n1583_ | ~new_n1587_ | ~new_n1591_ | ~new_n1595_;
  assign new_n1597_ = ~pi09 & ~pi10 & ~pi07;
  assign new_n1598_ = ~new_n1597_ | ~pi15 | ~new_n62_ | ~pi13;
  assign new_n1599_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1600_ = ~new_n24_ | ~pi02;
  assign new_n1601_ = ~new_n1600_ & ~pi03 & ~new_n1598_ & ~new_n1599_;
  assign new_n1602_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n1603_ = ~pi15 | ~new_n1602_ | ~pi13;
  assign new_n1604_ = ~pi02 | ~new_n66_ | ~new_n24_;
  assign new_n1605_ = ~new_n56_ & ~pi06 & ~new_n1603_ & ~new_n1604_;
  assign new_n1606_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n1607_ = ~pi15 | ~new_n1606_ | ~pi13;
  assign new_n1608_ = ~pi00 | ~new_n66_ | ~pi02;
  assign new_n1609_ = ~new_n56_ & ~pi06 & ~new_n1607_ & ~new_n1608_;
  assign new_n1610_ = ~new_n1609_ & ~new_n1605_ & ~new_n1596_ & ~new_n1601_;
  assign new_n1611_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1612_ = ~pi15 | ~new_n1611_ | ~pi13;
  assign new_n1613_ = ~pi00 | ~new_n66_ | ~pi02;
  assign new_n1614_ = ~new_n56_ & ~new_n64_ & ~new_n1612_ & ~new_n1613_;
  assign new_n1615_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n1616_ = ~pi15 | ~new_n1615_ | ~pi13;
  assign new_n1617_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1618_ = ~new_n56_ & ~new_n64_ & ~new_n1616_ & ~new_n1617_;
  assign new_n1619_ = ~pi09 & ~pi10 & ~pi07;
  assign new_n1620_ = ~new_n1619_ | ~pi15 | ~new_n62_ | ~pi13;
  assign new_n1621_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1622_ = ~new_n41_ | ~pi01;
  assign new_n1623_ = ~new_n1622_ & ~pi02 & ~new_n1620_ & ~new_n1621_;
  assign new_n1624_ = ~pi09 & ~pi10 & ~pi07;
  assign new_n1625_ = ~new_n1624_ | ~pi15 | ~new_n62_ | ~pi13;
  assign new_n1626_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1627_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1628_ = ~new_n1627_ & ~new_n1625_ & ~new_n1626_;
  assign new_n1629_ = ~new_n1628_ & ~new_n1623_ & ~new_n1614_ & ~new_n1618_;
  assign new_n1630_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n1631_ = ~pi15 | ~new_n1630_ | ~pi13;
  assign new_n1632_ = ~pi01 | ~new_n25_ | ~new_n41_;
  assign new_n1633_ = ~pi06 & ~pi05 & ~new_n1631_ & ~new_n1632_;
  assign new_n1634_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n1635_ = ~pi15 | ~new_n1634_ | ~pi13;
  assign new_n1636_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1637_ = ~pi06 & ~pi05 & ~new_n1635_ & ~new_n1636_;
  assign new_n1638_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n1639_ = ~pi15 | ~new_n1638_ | ~pi13;
  assign new_n1640_ = ~pi01 | ~new_n25_ | ~new_n41_;
  assign new_n1641_ = ~new_n56_ & ~pi06 & ~new_n1639_ & ~new_n1640_;
  assign new_n1642_ = ~pi10 & ~pi12 & ~pi09;
  assign new_n1643_ = ~pi15 | ~new_n1642_ | ~pi13;
  assign new_n1644_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1645_ = ~new_n56_ & ~pi06 & ~new_n1643_ & ~new_n1644_;
  assign new_n1646_ = ~new_n1645_ & ~new_n1641_ & ~new_n1633_ & ~new_n1637_;
  assign new_n1647_ = ~new_n1579_ | ~new_n1610_ | ~new_n1629_ | ~new_n1646_;
  assign new_n1648_ = ~pi06 & ~new_n56_;
  assign new_n1649_ = ~new_n1648_ | ~new_n66_ | ~pi02 | ~pi00;
  assign new_n1650_ = ~pi11 | ~new_n62_ | ~pi08;
  assign new_n1651_ = ~new_n26_ & ~pi14 & ~new_n1649_ & ~new_n1650_;
  assign new_n1652_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1653_ = ~new_n1652_ | ~pi06 | ~new_n56_ | ~pi05;
  assign new_n1654_ = ~new_n26_ & ~pi14 & ~pi12;
  assign new_n1655_ = ~new_n1654_ | ~pi11 | ~new_n64_ | ~pi08;
  assign new_n1656_ = ~new_n1653_ & ~new_n1655_;
  assign new_n1657_ = ~new_n26_ & ~pi14 & ~pi12;
  assign new_n1658_ = ~new_n1657_ | ~pi11 | ~new_n64_ | ~pi08;
  assign new_n1659_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1660_ = ~pi02 | ~pi00;
  assign new_n1661_ = ~new_n1660_ & ~pi03 & ~new_n1658_ & ~new_n1659_;
  assign new_n1662_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1663_ = ~pi07 | ~new_n1662_ | ~new_n104_;
  assign new_n1664_ = ~pi11 | ~new_n62_ | ~pi08;
  assign new_n1665_ = ~new_n26_ & ~pi14 & ~new_n1663_ & ~new_n1664_;
  assign new_n1666_ = ~new_n1665_ & ~new_n1661_ & ~new_n1651_ & ~new_n1656_;
  assign new_n1667_ = ~pi08 | ~pi11;
  assign new_n1668_ = ~new_n26_ & ~pi14 & ~pi12 & ~new_n1667_;
  assign new_n1669_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1670_ = ~new_n1668_ | ~new_n1669_ | ~pi07 | ~pi04;
  assign new_n1671_ = ~pi08 | ~pi11;
  assign new_n1672_ = ~new_n26_ & ~pi14 & ~pi12 & ~new_n1671_;
  assign new_n1673_ = ~new_n41_ & ~pi03 & ~new_n25_;
  assign new_n1674_ = ~new_n1672_ | ~new_n1673_ | ~new_n104_ | ~pi07;
  assign new_n1675_ = ~pi07 | ~pi04;
  assign new_n1676_ = ~new_n24_ & ~pi00 & ~new_n1675_ & ~pi02;
  assign new_n1677_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1678_ = ~new_n1676_ | ~new_n1677_ | ~new_n27_ | ~pi13;
  assign new_n1679_ = ~new_n1666_ | ~new_n1670_ | ~new_n1674_ | ~new_n1678_;
  assign new_n1680_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1681_ = ~pi06 & ~new_n1680_ & ~pi05;
  assign new_n1682_ = ~new_n22_ & ~pi12 & ~new_n89_;
  assign new_n1683_ = ~new_n1681_ | ~new_n1682_ | ~new_n27_ | ~pi13;
  assign new_n1684_ = ~pi08 | ~pi11;
  assign new_n1685_ = ~new_n26_ & ~pi14 & ~pi12 & ~new_n1684_;
  assign new_n1686_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1687_ = ~new_n1685_ | ~new_n1686_ | ~new_n57_ | ~pi04;
  assign new_n1688_ = ~pi08 | ~pi11;
  assign new_n1689_ = ~new_n26_ & ~pi14 & ~pi12 & ~new_n1688_;
  assign new_n1690_ = ~new_n24_ & ~new_n66_ & ~pi00;
  assign new_n1691_ = ~new_n1689_ | ~new_n1690_ | ~new_n57_ | ~pi04;
  assign new_n1692_ = ~pi08 | ~pi11;
  assign new_n1693_ = ~new_n26_ & ~pi14 & ~pi12 & ~new_n1692_;
  assign new_n1694_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1695_ = ~new_n1693_ | ~new_n1694_ | ~new_n104_ | ~pi07;
  assign new_n1696_ = ~new_n1683_ | ~new_n1687_ | ~new_n1691_ | ~new_n1695_;
  assign new_n1697_ = ~pi08 | ~pi11;
  assign new_n1698_ = ~new_n26_ & ~pi14 & ~pi12 & ~new_n1697_;
  assign new_n1699_ = ~new_n24_ & ~new_n66_ & ~pi00;
  assign new_n1700_ = ~new_n1698_ | ~new_n1699_ | ~new_n104_ | ~pi07;
  assign new_n1701_ = ~pi08 | ~pi11;
  assign new_n1702_ = ~new_n26_ & ~pi14 & ~pi12 & ~new_n1701_;
  assign new_n1703_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1704_ = ~new_n1702_ | ~new_n1703_ | ~new_n104_ | ~new_n57_;
  assign new_n1705_ = ~pi02 | ~pi00;
  assign new_n1706_ = ~pi06 & ~pi05 & ~pi03 & ~new_n1705_;
  assign new_n1707_ = ~new_n22_ & ~pi12 & ~new_n89_;
  assign new_n1708_ = ~new_n1706_ | ~new_n1707_ | ~new_n27_ | ~pi13;
  assign new_n1709_ = ~pi08 | ~pi11;
  assign new_n1710_ = ~new_n26_ & ~pi14 & ~pi12 & ~new_n1709_;
  assign new_n1711_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1712_ = ~new_n1710_ | ~new_n1711_ | ~new_n57_ | ~pi04;
  assign new_n1713_ = ~new_n1700_ | ~new_n1704_ | ~new_n1708_ | ~new_n1712_;
  assign new_n1714_ = ~new_n1713_ & ~new_n1679_ & ~new_n1696_;
  assign new_n1715_ = ~pi13 | ~pi15;
  assign new_n1716_ = ~new_n22_ & ~pi09 & ~new_n1715_ & ~pi12;
  assign new_n1717_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1718_ = ~new_n1716_ | ~new_n1717_ | ~pi07 | ~pi04;
  assign new_n1719_ = ~pi13 | ~pi15;
  assign new_n1720_ = ~new_n22_ & ~pi09 & ~new_n1719_ & ~pi12;
  assign new_n1721_ = ~new_n41_ & ~pi03 & ~new_n25_;
  assign new_n1722_ = ~new_n1720_ | ~new_n1721_ | ~pi07 | ~pi04;
  assign new_n1723_ = ~pi08 | ~pi11;
  assign new_n1724_ = ~new_n26_ & ~pi14 & ~pi12 & ~new_n1723_;
  assign new_n1725_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1726_ = ~new_n1724_ | ~new_n1725_ | ~pi07 | ~pi04;
  assign new_n1727_ = ~pi08 | ~pi11;
  assign new_n1728_ = ~new_n26_ & ~pi14 & ~pi12 & ~new_n1727_;
  assign new_n1729_ = ~new_n24_ & ~new_n66_ & ~pi00;
  assign new_n1730_ = ~new_n1728_ | ~new_n1729_ | ~pi07 | ~pi04;
  assign new_n1731_ = ~new_n1718_ | ~new_n1722_ | ~new_n1726_ | ~new_n1730_;
  assign new_n1732_ = ~pi05 & ~pi06;
  assign new_n1733_ = ~new_n1732_ | ~new_n25_ | ~new_n41_ | ~pi01;
  assign new_n1734_ = ~pi11 | ~new_n62_ | ~pi08;
  assign new_n1735_ = ~new_n26_ & ~pi14 & ~new_n1733_ & ~new_n1734_;
  assign new_n1736_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1737_ = ~new_n1736_ | ~pi06 | ~new_n56_ | ~pi05;
  assign new_n1738_ = ~new_n26_ & ~pi14 & ~pi12;
  assign new_n1739_ = ~new_n1738_ | ~pi11 | ~new_n64_ | ~pi08;
  assign new_n1740_ = ~new_n1737_ & ~new_n1739_;
  assign new_n1741_ = ~new_n26_ & ~pi14 & ~pi12;
  assign new_n1742_ = ~new_n1741_ | ~pi11 | ~new_n64_ | ~pi08;
  assign new_n1743_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1744_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1745_ = ~new_n1744_ & ~new_n1742_ & ~new_n1743_;
  assign new_n1746_ = ~new_n1745_ & ~new_n1740_ & ~new_n1731_ & ~new_n1735_;
  assign new_n1747_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1748_ = ~pi15 | ~new_n1747_ | ~pi13;
  assign new_n1749_ = ~pi02 | ~new_n66_ | ~new_n24_;
  assign new_n1750_ = ~pi06 & ~pi05 & ~new_n1748_ & ~new_n1749_;
  assign new_n1751_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1752_ = ~pi15 | ~new_n1751_ | ~pi13;
  assign new_n1753_ = ~pi00 | ~new_n66_ | ~pi02;
  assign new_n1754_ = ~pi06 & ~pi05 & ~new_n1752_ & ~new_n1753_;
  assign new_n1755_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1756_ = ~pi15 | ~new_n1755_ | ~pi13;
  assign new_n1757_ = ~pi02 | ~new_n66_ | ~new_n24_;
  assign new_n1758_ = ~new_n56_ & ~pi06 & ~new_n1756_ & ~new_n1757_;
  assign new_n1759_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1760_ = ~pi15 | ~new_n1759_ | ~pi13;
  assign new_n1761_ = ~pi00 | ~new_n66_ | ~pi02;
  assign new_n1762_ = ~new_n56_ & ~pi06 & ~new_n1760_ & ~new_n1761_;
  assign new_n1763_ = ~new_n1762_ & ~new_n1758_ & ~new_n1750_ & ~new_n1754_;
  assign new_n1764_ = ~pi09 & ~new_n22_ & ~pi07;
  assign new_n1765_ = ~new_n1764_ | ~pi15 | ~new_n62_ | ~pi13;
  assign new_n1766_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1767_ = ~new_n24_ | ~pi02;
  assign new_n1768_ = ~new_n1767_ & ~pi03 & ~new_n1765_ & ~new_n1766_;
  assign new_n1769_ = ~pi09 & ~new_n22_ & ~pi07;
  assign new_n1770_ = ~new_n1769_ | ~pi15 | ~new_n62_ | ~pi13;
  assign new_n1771_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1772_ = ~pi02 | ~pi00;
  assign new_n1773_ = ~new_n1772_ & ~pi03 & ~new_n1770_ & ~new_n1771_;
  assign new_n1774_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1775_ = ~pi15 | ~new_n1774_ | ~pi13;
  assign new_n1776_ = ~pi02 | ~new_n66_ | ~new_n24_;
  assign new_n1777_ = ~new_n64_ & ~pi05 & ~new_n1775_ & ~new_n1776_;
  assign new_n1778_ = ~new_n22_ & ~pi12 & ~pi09;
  assign new_n1779_ = ~pi15 | ~new_n1778_ | ~pi13;
  assign new_n1780_ = ~pi00 | ~new_n66_ | ~pi02;
  assign new_n1781_ = ~new_n64_ & ~pi05 & ~new_n1779_ & ~new_n1780_;
  assign new_n1782_ = ~new_n1781_ & ~new_n1777_ & ~new_n1768_ & ~new_n1773_;
  assign new_n1783_ = ~new_n1714_ | ~new_n1746_ | ~new_n1763_ | ~new_n1782_;
  assign new_n1784_ = ~pi08 | ~pi11;
  assign new_n1785_ = ~new_n26_ & ~pi14 & ~pi12 & ~new_n1784_;
  assign new_n1786_ = ~new_n41_ & ~pi03 & ~new_n25_;
  assign new_n1787_ = ~new_n1785_ | ~new_n1786_ | ~pi07 | ~pi04;
  assign new_n1788_ = ~pi07 | ~pi04;
  assign new_n1789_ = ~new_n24_ & ~pi00 & ~new_n1788_ & ~new_n66_;
  assign new_n1790_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1791_ = ~new_n1789_ | ~new_n1790_ | ~new_n27_ | ~pi13;
  assign new_n1792_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1793_ = ~new_n24_ & ~pi00 & ~new_n1792_ & ~pi02;
  assign new_n1794_ = ~new_n89_ & ~pi10 & ~pi07;
  assign new_n1795_ = ~new_n26_ & ~pi14 & ~pi12;
  assign new_n1796_ = ~new_n1795_ | ~new_n1793_ | ~new_n1794_;
  assign new_n1797_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1798_ = ~new_n24_ & ~pi00 & ~new_n1797_ & ~new_n66_;
  assign new_n1799_ = ~new_n89_ & ~pi10 & ~pi07;
  assign new_n1800_ = ~new_n26_ & ~pi14 & ~pi12;
  assign new_n1801_ = ~new_n1800_ | ~new_n1798_ | ~new_n1799_;
  assign new_n1802_ = ~new_n1787_ | ~new_n1791_ | ~new_n1796_ | ~new_n1801_;
  assign new_n1803_ = ~new_n41_ | ~pi01;
  assign new_n1804_ = ~pi06 & ~pi05 & ~pi02 & ~new_n1803_;
  assign new_n1805_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1806_ = ~new_n1804_ | ~new_n1805_ | ~new_n27_ | ~pi13;
  assign new_n1807_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1808_ = ~pi06 & ~new_n1807_ & ~pi05;
  assign new_n1809_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1810_ = ~new_n1808_ | ~new_n1809_ | ~new_n27_ | ~pi13;
  assign new_n1811_ = ~new_n57_ | ~pi04;
  assign new_n1812_ = ~new_n24_ & ~pi00 & ~new_n1811_ & ~pi02;
  assign new_n1813_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1814_ = ~new_n1812_ | ~new_n1813_ | ~new_n27_ | ~pi13;
  assign new_n1815_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1816_ = ~new_n56_ & ~new_n1815_ & ~pi06;
  assign new_n1817_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1818_ = ~new_n1816_ | ~new_n1817_ | ~new_n27_ | ~pi13;
  assign new_n1819_ = ~new_n1806_ | ~new_n1810_ | ~new_n1814_ | ~new_n1818_;
  assign new_n1820_ = ~new_n104_ | ~pi07;
  assign new_n1821_ = ~new_n24_ & ~pi00 & ~new_n1820_ & ~pi02;
  assign new_n1822_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1823_ = ~new_n1821_ | ~new_n1822_ | ~new_n27_ | ~pi13;
  assign new_n1824_ = ~pi01 | ~pi03 | ~new_n41_;
  assign new_n1825_ = ~new_n64_ & ~new_n1824_ & ~pi05;
  assign new_n1826_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1827_ = ~new_n1825_ | ~new_n1826_ | ~new_n27_ | ~pi13;
  assign new_n1828_ = ~new_n24_ | ~pi02;
  assign new_n1829_ = ~pi06 & ~pi05 & ~pi03 & ~new_n1828_;
  assign new_n1830_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1831_ = ~new_n1829_ | ~new_n1830_ | ~new_n27_ | ~pi13;
  assign new_n1832_ = ~pi02 | ~pi00;
  assign new_n1833_ = ~pi06 & ~pi05 & ~pi03 & ~new_n1832_;
  assign new_n1834_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1835_ = ~new_n1833_ | ~new_n1834_ | ~new_n27_ | ~pi13;
  assign new_n1836_ = ~new_n1823_ | ~new_n1827_ | ~new_n1831_ | ~new_n1835_;
  assign new_n1837_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1838_ = ~new_n25_ & ~pi01 & ~new_n1837_ & ~pi03;
  assign new_n1839_ = ~new_n89_ & ~pi10 & ~pi07;
  assign new_n1840_ = ~new_n26_ & ~pi14 & ~pi12;
  assign new_n1841_ = ~new_n1840_ | ~new_n1838_ | ~new_n1839_;
  assign new_n1842_ = ~new_n57_ | ~pi04;
  assign new_n1843_ = ~new_n25_ & ~pi01 & ~new_n1842_ & ~pi03;
  assign new_n1844_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1845_ = ~new_n1843_ | ~new_n1844_ | ~new_n27_ | ~pi13;
  assign new_n1846_ = ~pi02 | ~pi00;
  assign new_n1847_ = ~new_n56_ & ~pi06 & ~pi03 & ~new_n1846_;
  assign new_n1848_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1849_ = ~new_n1847_ | ~new_n1848_ | ~new_n27_ | ~pi13;
  assign new_n1850_ = ~new_n1849_ | ~new_n1841_ | ~new_n1845_;
  assign new_n1851_ = ~new_n1850_ & ~new_n1836_ & ~new_n1802_ & ~new_n1819_;
  assign new_n1852_ = ~new_n41_ | ~pi01 | ~new_n56_ | ~pi03;
  assign new_n1853_ = ~new_n104_ & ~new_n57_ & ~new_n1852_ & ~pi07;
  assign new_n1854_ = ~new_n19_ & ~pi11 & ~pi08 & ~new_n79_;
  assign new_n1855_ = ~pi12 & ~new_n26_;
  assign new_n1856_ = ~new_n1853_ | ~new_n1854_ | ~pi15 | ~new_n1855_;
  assign new_n1857_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1858_ = ~new_n26_ & ~pi12 & ~new_n1857_ & ~new_n37_;
  assign new_n1859_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1860_ = ~pi06 & ~pi08 & ~pi05;
  assign new_n1861_ = ~new_n1860_ | ~new_n1858_ | ~new_n1859_;
  assign new_n1862_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1863_ = ~new_n26_ & ~pi12 & ~new_n1862_ & ~new_n37_;
  assign new_n1864_ = ~pi06 & ~pi08 & ~pi05;
  assign new_n1865_ = ~pi00 & ~new_n24_;
  assign new_n1866_ = ~new_n1863_ | ~new_n1864_ | ~pi03 | ~new_n1865_;
  assign new_n1867_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1868_ = ~new_n26_ & ~pi12 & ~new_n1867_ & ~new_n37_;
  assign new_n1869_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1870_ = ~new_n56_ & ~pi08 & ~pi06;
  assign new_n1871_ = ~new_n1870_ | ~new_n1868_ | ~new_n1869_;
  assign new_n1872_ = ~new_n1856_ | ~new_n1861_ | ~new_n1866_ | ~new_n1871_;
  assign new_n1873_ = ~new_n64_ & ~pi08 & ~pi05;
  assign new_n1874_ = ~new_n1873_ | ~pi03 | ~new_n41_ | ~pi01;
  assign new_n1875_ = ~pi13 | ~pi15 | ~new_n62_;
  assign new_n1876_ = ~pi09 | ~pi10;
  assign new_n1877_ = ~new_n1876_ & ~pi11 & ~new_n1874_ & ~new_n1875_;
  assign new_n1878_ = ~new_n56_ & ~pi08 & ~pi06;
  assign new_n1879_ = ~new_n1878_ | ~pi03 | ~new_n41_ | ~pi01;
  assign new_n1880_ = ~pi13 | ~pi15 | ~new_n62_;
  assign new_n1881_ = ~pi09 | ~pi10;
  assign new_n1882_ = ~new_n1881_ & ~pi11 & ~new_n1879_ & ~new_n1880_;
  assign new_n1883_ = ~new_n64_ & ~pi08 & ~pi05;
  assign new_n1884_ = ~new_n1883_ | ~new_n25_ | ~new_n41_ | ~pi01;
  assign new_n1885_ = ~pi13 | ~pi15 | ~new_n62_;
  assign new_n1886_ = ~pi09 | ~pi10;
  assign new_n1887_ = ~new_n1886_ & ~pi11 & ~new_n1884_ & ~new_n1885_;
  assign new_n1888_ = ~new_n1887_ & ~new_n1882_ & ~new_n1872_ & ~new_n1877_;
  assign new_n1889_ = ~new_n89_ & ~pi10 & ~pi07;
  assign new_n1890_ = ~new_n1889_ | ~new_n27_ | ~new_n62_ | ~pi13;
  assign new_n1891_ = ~pi05 | ~pi06 | ~new_n56_;
  assign new_n1892_ = ~pi02 | ~pi00;
  assign new_n1893_ = ~new_n1892_ & ~pi03 & ~new_n1890_ & ~new_n1891_;
  assign new_n1894_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1895_ = ~pi13 | ~new_n1894_ | ~new_n27_;
  assign new_n1896_ = ~pi02 | ~new_n66_ | ~new_n24_;
  assign new_n1897_ = ~new_n64_ & ~pi05 & ~new_n1895_ & ~new_n1896_;
  assign new_n1898_ = ~new_n89_ & ~pi12 & ~pi10;
  assign new_n1899_ = ~pi13 | ~new_n1898_ | ~new_n27_;
  assign new_n1900_ = ~pi00 | ~new_n66_ | ~pi02;
  assign new_n1901_ = ~new_n64_ & ~pi05 & ~new_n1899_ & ~new_n1900_;
  assign new_n1902_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1903_ = ~pi04 | ~new_n1902_ | ~pi07;
  assign new_n1904_ = ~pi08 | ~new_n62_ | ~new_n19_;
  assign new_n1905_ = ~new_n26_ & ~pi14 & ~new_n1903_ & ~new_n1904_;
  assign new_n1906_ = ~new_n1905_ & ~new_n1901_ & ~new_n1893_ & ~new_n1897_;
  assign new_n1907_ = ~new_n41_ & ~pi03 & ~new_n25_;
  assign new_n1908_ = ~pi04 | ~new_n1907_ | ~pi07;
  assign new_n1909_ = ~pi08 | ~new_n62_ | ~new_n19_;
  assign new_n1910_ = ~new_n26_ & ~pi14 & ~new_n1908_ & ~new_n1909_;
  assign new_n1911_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1912_ = ~new_n1911_ | ~new_n89_ | ~pi07 | ~pi04;
  assign new_n1913_ = ~pi13 | ~pi15 | ~new_n62_;
  assign new_n1914_ = ~pi09 | ~pi10;
  assign new_n1915_ = ~new_n1914_ & ~pi11 & ~new_n1912_ & ~new_n1913_;
  assign new_n1916_ = ~new_n24_ & ~new_n66_ & ~pi00;
  assign new_n1917_ = ~new_n1916_ | ~new_n89_ | ~pi07 | ~pi04;
  assign new_n1918_ = ~pi13 | ~pi15 | ~new_n62_;
  assign new_n1919_ = ~pi09 | ~pi10;
  assign new_n1920_ = ~new_n1919_ & ~pi11 & ~new_n1917_ & ~new_n1918_;
  assign new_n1921_ = ~pi04 & ~pi02 & ~pi00 & ~new_n24_;
  assign new_n1922_ = ~new_n1921_ | ~new_n64_ | ~pi06 | ~pi05;
  assign new_n1923_ = ~new_n19_ & ~pi11 & ~pi08 & ~new_n79_;
  assign new_n1924_ = ~new_n1923_ | ~pi15 | ~new_n62_ | ~pi13;
  assign new_n1925_ = ~new_n1922_ & ~new_n1924_;
  assign new_n1926_ = ~new_n1925_ & ~new_n1920_ & ~new_n1910_ & ~new_n1915_;
  assign new_n1927_ = ~new_n1851_ | ~new_n1888_ | ~new_n1906_ | ~new_n1926_;
  assign new_n1928_ = ~new_n56_ & ~pi08 & ~pi06;
  assign new_n1929_ = ~new_n1928_ | ~new_n66_ | ~pi02 | ~pi00;
  assign new_n1930_ = ~pi13 | ~new_n27_ | ~new_n62_;
  assign new_n1931_ = ~pi09 | ~pi10;
  assign new_n1932_ = ~new_n1931_ & ~pi11 & ~new_n1929_ & ~new_n1930_;
  assign new_n1933_ = ~pi04 & ~pi03 & ~pi01 & ~new_n25_;
  assign new_n1934_ = ~new_n1933_ | ~new_n64_ | ~pi06 | ~pi05;
  assign new_n1935_ = ~new_n89_ | ~pi09 | ~new_n22_ | ~pi10;
  assign new_n1936_ = ~new_n62_ | ~pi13;
  assign new_n1937_ = ~new_n1936_ & ~pi14 & ~new_n1934_ & ~new_n1935_;
  assign new_n1938_ = ~new_n19_ & ~pi11 & ~pi08 & ~new_n79_;
  assign new_n1939_ = ~new_n1938_ | ~new_n27_ | ~new_n62_ | ~pi13;
  assign new_n1940_ = ~pi02 | ~pi00 | ~new_n66_ | ~new_n56_;
  assign new_n1941_ = ~pi06 | ~pi05;
  assign new_n1942_ = ~new_n1941_ & ~pi07 & ~new_n1939_ & ~new_n1940_;
  assign new_n1943_ = ~new_n64_ & ~pi08 & ~pi05;
  assign new_n1944_ = ~new_n1943_ | ~new_n66_ | ~new_n24_ | ~pi02;
  assign new_n1945_ = ~pi13 | ~new_n27_ | ~new_n62_;
  assign new_n1946_ = ~pi09 | ~pi10;
  assign new_n1947_ = ~new_n1946_ & ~pi11 & ~new_n1944_ & ~new_n1945_;
  assign new_n1948_ = ~new_n1947_ & ~new_n1942_ & ~new_n1932_ & ~new_n1937_;
  assign new_n1949_ = ~pi04 | ~new_n89_ | ~pi07;
  assign new_n1950_ = ~new_n41_ & ~new_n25_ & ~new_n1949_ & ~pi03;
  assign new_n1951_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1952_ = ~new_n26_ & ~pi12 & ~new_n1951_ & ~pi14;
  assign new_n1953_ = ~new_n1950_ | ~new_n1952_;
  assign new_n1954_ = ~pi00 | ~new_n66_ | ~pi02;
  assign new_n1955_ = ~new_n64_ & ~pi05 & ~new_n1954_ & ~pi08;
  assign new_n1956_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1957_ = ~new_n26_ & ~pi12 & ~new_n1956_ & ~pi14;
  assign new_n1958_ = ~new_n1955_ | ~new_n1957_;
  assign new_n1959_ = ~pi04 | ~new_n89_ | ~pi07;
  assign new_n1960_ = ~new_n25_ & ~pi01 & ~new_n1959_ & ~pi03;
  assign new_n1961_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1962_ = ~new_n26_ & ~pi12 & ~new_n1961_ & ~pi14;
  assign new_n1963_ = ~new_n1960_ | ~new_n1962_;
  assign new_n1964_ = ~new_n1948_ | ~new_n1953_ | ~new_n1958_ | ~new_n1963_;
  assign new_n1965_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1966_ = ~new_n26_ & ~pi12 & ~new_n1965_ & ~pi14;
  assign new_n1967_ = ~pi06 & ~pi08 & ~pi05;
  assign new_n1968_ = ~pi00 & ~new_n24_;
  assign new_n1969_ = ~new_n1966_ | ~new_n1967_ | ~pi03 | ~new_n1968_;
  assign new_n1970_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1971_ = ~new_n26_ & ~pi12 & ~new_n1970_ & ~pi14;
  assign new_n1972_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1973_ = ~new_n56_ & ~pi08 & ~pi06;
  assign new_n1974_ = ~new_n1973_ | ~new_n1971_ | ~new_n1972_;
  assign new_n1975_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1976_ = ~new_n26_ & ~pi12 & ~new_n1975_ & ~pi14;
  assign new_n1977_ = ~new_n56_ & ~pi08 & ~pi06;
  assign new_n1978_ = ~pi00 & ~new_n24_;
  assign new_n1979_ = ~new_n1976_ | ~new_n1977_ | ~pi03 | ~new_n1978_;
  assign new_n1980_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1981_ = ~new_n26_ & ~pi12 & ~new_n1980_ & ~pi14;
  assign new_n1982_ = ~new_n24_ & ~pi02 & ~pi00;
  assign new_n1983_ = ~new_n64_ & ~pi08 & ~pi05;
  assign new_n1984_ = ~new_n1983_ | ~new_n1981_ | ~new_n1982_;
  assign new_n1985_ = ~new_n1969_ | ~new_n1974_ | ~new_n1979_ | ~new_n1984_;
  assign new_n1986_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1987_ = ~new_n26_ & ~pi12 & ~new_n1986_ & ~pi14;
  assign new_n1988_ = ~new_n64_ & ~pi08 & ~pi05;
  assign new_n1989_ = ~pi00 & ~new_n24_;
  assign new_n1990_ = ~new_n1987_ | ~new_n1988_ | ~pi03 | ~new_n1989_;
  assign new_n1991_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1992_ = ~new_n26_ & ~pi12 & ~new_n1991_ & ~pi14;
  assign new_n1993_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n1994_ = ~pi06 & ~pi08 & ~pi05;
  assign new_n1995_ = ~new_n1994_ | ~new_n1992_ | ~new_n1993_;
  assign new_n1996_ = ~pi00 | ~new_n66_ | ~pi02;
  assign new_n1997_ = ~pi06 & ~pi05 & ~new_n1996_ & ~pi08;
  assign new_n1998_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n1999_ = ~new_n26_ & ~pi12 & ~new_n1998_ & ~pi14;
  assign new_n2000_ = ~new_n1997_ | ~new_n1999_;
  assign new_n2001_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n2002_ = ~new_n26_ & ~pi12 & ~new_n2001_ & ~pi14;
  assign new_n2003_ = ~new_n25_ & ~pi03 & ~pi01;
  assign new_n2004_ = ~new_n56_ & ~pi08 & ~pi06;
  assign new_n2005_ = ~new_n2004_ | ~new_n2002_ | ~new_n2003_;
  assign new_n2006_ = ~new_n1990_ | ~new_n1995_ | ~new_n2000_ | ~new_n2005_;
  assign new_n2007_ = ~new_n2006_ & ~new_n1964_ & ~new_n1985_;
  assign new_n2008_ = ~pi04 | ~new_n89_ | ~pi07;
  assign new_n2009_ = ~new_n24_ & ~pi00 & ~new_n2008_ & ~pi02;
  assign new_n2010_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n2011_ = ~new_n26_ & ~pi12 & ~new_n2010_ & ~pi14;
  assign new_n2012_ = ~new_n2009_ | ~new_n2011_;
  assign new_n2013_ = ~pi04 | ~new_n89_ | ~pi07;
  assign new_n2014_ = ~new_n25_ & ~pi01 & ~new_n2013_ & ~pi03;
  assign new_n2015_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n2016_ = ~new_n26_ & ~pi12 & ~new_n2015_ & ~new_n37_;
  assign new_n2017_ = ~new_n2014_ | ~new_n2016_;
  assign new_n2018_ = ~pi04 | ~new_n89_ | ~pi07;
  assign new_n2019_ = ~new_n41_ & ~new_n25_ & ~new_n2018_ & ~pi03;
  assign new_n2020_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n2021_ = ~new_n26_ & ~pi12 & ~new_n2020_ & ~new_n37_;
  assign new_n2022_ = ~new_n2019_ | ~new_n2021_;
  assign new_n2023_ = ~pi04 | ~new_n89_ | ~pi07;
  assign new_n2024_ = ~new_n24_ & ~pi00 & ~new_n2023_ & ~new_n66_;
  assign new_n2025_ = ~pi10 | ~new_n22_ | ~pi09;
  assign new_n2026_ = ~new_n26_ & ~pi12 & ~new_n2025_ & ~pi14;
  assign new_n2027_ = ~new_n2024_ | ~new_n2026_;
  assign new_n2028_ = ~new_n2012_ | ~new_n2017_ | ~new_n2022_ | ~new_n2027_;
  assign new_n2029_ = ~pi06 & ~pi08 & ~pi05;
  assign new_n2030_ = ~new_n2029_ | ~new_n25_ | ~new_n41_ | ~pi01;
  assign new_n2031_ = ~pi13 | ~new_n27_ | ~new_n62_;
  assign new_n2032_ = ~pi09 | ~pi10;
  assign new_n2033_ = ~new_n2032_ & ~pi11 & ~new_n2030_ & ~new_n2031_;
  assign new_n2034_ = ~pi04 & ~pi02 & ~pi00 & ~new_n24_;
  assign new_n2035_ = ~new_n2034_ | ~new_n64_ | ~pi06 | ~pi05;
  assign new_n2036_ = ~new_n89_ | ~pi09 | ~new_n22_ | ~pi10;
  assign new_n2037_ = ~new_n62_ | ~pi13;
  assign new_n2038_ = ~new_n2037_ & ~pi14 & ~new_n2035_ & ~new_n2036_;
  assign new_n2039_ = ~new_n19_ & ~pi11 & ~pi08 & ~new_n79_;
  assign new_n2040_ = ~new_n2039_ | ~new_n27_ | ~new_n62_ | ~pi13;
  assign new_n2041_ = ~new_n41_ | ~pi01 | ~new_n56_ | ~pi03;
  assign new_n2042_ = ~pi06 | ~pi05;
  assign new_n2043_ = ~new_n2042_ & ~pi07 & ~new_n2040_ & ~new_n2041_;
  assign new_n2044_ = ~new_n2043_ & ~new_n2038_ & ~new_n2028_ & ~new_n2033_;
  assign new_n2045_ = ~pi06 & ~pi08 & ~pi05;
  assign new_n2046_ = ~new_n2045_ | ~new_n66_ | ~new_n24_ | ~pi02;
  assign new_n2047_ = ~pi13 | ~pi15 | ~new_n62_;
  assign new_n2048_ = ~pi09 | ~pi10;
  assign new_n2049_ = ~new_n2048_ & ~pi11 & ~new_n2046_ & ~new_n2047_;
  assign new_n2050_ = ~pi06 & ~pi08 & ~pi05;
  assign new_n2051_ = ~new_n2050_ | ~new_n66_ | ~pi02 | ~pi00;
  assign new_n2052_ = ~pi13 | ~pi15 | ~new_n62_;
  assign new_n2053_ = ~pi09 | ~pi10;
  assign new_n2054_ = ~new_n2053_ & ~pi11 & ~new_n2051_ & ~new_n2052_;
  assign new_n2055_ = ~new_n56_ & ~pi08 & ~pi06;
  assign new_n2056_ = ~new_n2055_ | ~new_n66_ | ~new_n24_ | ~pi02;
  assign new_n2057_ = ~pi13 | ~pi15 | ~new_n62_;
  assign new_n2058_ = ~pi09 | ~pi10;
  assign new_n2059_ = ~new_n2058_ & ~pi11 & ~new_n2056_ & ~new_n2057_;
  assign new_n2060_ = ~new_n56_ & ~pi08 & ~pi06;
  assign new_n2061_ = ~new_n2060_ | ~new_n66_ | ~pi02 | ~pi00;
  assign new_n2062_ = ~pi13 | ~pi15 | ~new_n62_;
  assign new_n2063_ = ~pi09 | ~pi10;
  assign new_n2064_ = ~new_n2063_ & ~pi11 & ~new_n2061_ & ~new_n2062_;
  assign new_n2065_ = ~new_n2064_ & ~new_n2059_ & ~new_n2049_ & ~new_n2054_;
  assign new_n2066_ = ~pi04 & ~pi03 & ~pi01 & ~new_n25_;
  assign new_n2067_ = ~new_n2066_ | ~new_n64_ | ~pi06 | ~pi05;
  assign new_n2068_ = ~new_n19_ & ~pi11 & ~pi08 & ~new_n79_;
  assign new_n2069_ = ~new_n2068_ | ~pi15 | ~new_n62_ | ~pi13;
  assign new_n2070_ = ~new_n2067_ & ~new_n2069_;
  assign new_n2071_ = ~new_n19_ & ~pi11 & ~pi08 & ~new_n79_;
  assign new_n2072_ = ~new_n2071_ | ~pi15 | ~new_n62_ | ~pi13;
  assign new_n2073_ = ~pi02 | ~pi00 | ~new_n66_ | ~new_n56_;
  assign new_n2074_ = ~pi06 | ~pi05;
  assign new_n2075_ = ~new_n2074_ & ~pi07 & ~new_n2072_ & ~new_n2073_;
  assign new_n2076_ = ~new_n64_ & ~pi08 & ~pi05;
  assign new_n2077_ = ~new_n2076_ | ~new_n66_ | ~new_n24_ | ~pi02;
  assign new_n2078_ = ~pi13 | ~pi15 | ~new_n62_;
  assign new_n2079_ = ~pi09 | ~pi10;
  assign new_n2080_ = ~new_n2079_ & ~pi11 & ~new_n2077_ & ~new_n2078_;
  assign new_n2081_ = ~new_n64_ & ~pi08 & ~pi05;
  assign new_n2082_ = ~new_n2081_ | ~new_n66_ | ~pi02 | ~pi00;
  assign new_n2083_ = ~pi13 | ~pi15 | ~new_n62_;
  assign new_n2084_ = ~pi09 | ~pi10;
  assign new_n2085_ = ~new_n2084_ & ~pi11 & ~new_n2082_ & ~new_n2083_;
  assign new_n2086_ = ~new_n2085_ & ~new_n2080_ & ~new_n2070_ & ~new_n2075_;
  assign new_n2087_ = ~new_n2007_ | ~new_n2044_ | ~new_n2065_ | ~new_n2086_;
  assign new_n2088_ = ~new_n2087_ & ~new_n1927_ & ~new_n1647_ & ~new_n1783_;
  assign po0 = ~new_n389_ | ~new_n934_ | ~new_n1511_ | ~new_n2088_;
endmodule


