// Benchmark "i8" written by ABC on Thu Mar 19 13:02:36 2020

module i8 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47,
    po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71,
    po72, po73, po74, po75, po76, po77, po78, po79, po80  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46,
    po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58,
    po59, po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70,
    po71, po72, po73, po74, po75, po76, po77, po78, po79, po80;
  wire new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n571_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n596_,
    new_n598_, new_n600_, new_n602_, new_n604_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n663_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n721_, new_n723_, new_n725_, new_n727_, new_n729_,
    new_n731_, new_n733_, new_n735_, new_n737_, new_n739_, new_n741_,
    new_n743_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n862_, new_n864_, new_n866_, new_n868_,
    new_n870_, new_n872_, new_n874_, new_n876_, new_n878_, new_n880_,
    new_n882_, new_n884_, new_n886_, new_n888_, new_n890_, new_n892_,
    new_n894_, new_n896_, new_n898_, new_n900_, new_n902_, new_n904_,
    new_n906_, new_n908_, new_n910_, new_n912_, new_n914_, new_n916_,
    new_n918_, new_n920_, new_n922_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1107_,
    new_n1109_, new_n1111_, new_n1113_, new_n1115_, new_n1117_, new_n1119_,
    new_n1121_, new_n1123_, new_n1125_, new_n1127_, new_n1129_, new_n1131_,
    new_n1133_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_,
    new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_,
    new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_,
    new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_,
    new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_,
    new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_,
    new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_,
    new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_,
    new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_,
    new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_,
    new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_,
    new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_,
    new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_,
    new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_,
    new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_,
    new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_,
    new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_,
    new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_,
    new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_,
    new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_,
    new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_,
    new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_,
    new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_,
    new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_,
    new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_,
    new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_,
    new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_,
    new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_,
    new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_,
    new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_,
    new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_,
    new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_,
    new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_,
    new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_,
    new_n1394_, new_n1395_, new_n1396_, new_n1397_;
  assign new_n215_ = pi002 & pi000 & pi001;
  assign new_n216_ = ~pi003;
  assign new_n217_ = ~pi004;
  assign new_n218_ = ~pi005;
  assign new_n219_ = new_n217_ & new_n218_ & new_n216_;
  assign new_n220_ = ~pi002;
  assign new_n221_ = ~pi006;
  assign new_n222_ = new_n221_ & new_n220_ & pi001 & new_n218_ & new_n217_;
  assign new_n223_ = pi007 & new_n218_ & new_n216_;
  assign new_n224_ = pi008 & new_n218_ & pi001;
  assign new_n225_ = ~pi000;
  assign new_n226_ = new_n225_ & pi001 & new_n218_ & pi002;
  assign new_n227_ = ~pi001;
  assign new_n228_ = new_n221_ & pi002 & pi003 & new_n227_ & new_n218_ & new_n217_;
  assign new_n229_ = pi008 & new_n227_ & new_n218_ & pi002;
  assign new_n230_ = new_n221_ & new_n220_ & new_n227_ & new_n218_ & new_n217_;
  assign new_n231_ = pi007 & new_n227_ & new_n218_ & new_n220_;
  assign new_n232_ = pi005 | new_n215_;
  assign new_n233_ = new_n224_ | new_n222_ | new_n219_ | new_n223_;
  assign new_n234_ = new_n228_ | new_n229_ | new_n226_;
  assign new_n235_ = new_n231_ | new_n230_;
  assign new_n236_ = new_n232_ & pi009;
  assign new_n237_ = new_n232_ & pi010;
  assign new_n238_ = new_n232_ & pi011;
  assign new_n239_ = new_n232_ & pi012;
  assign new_n240_ = new_n232_ & pi013;
  assign new_n241_ = new_n232_ & pi014;
  assign new_n242_ = new_n232_ & pi015;
  assign new_n243_ = new_n232_ & pi016;
  assign new_n244_ = new_n232_ & pi017;
  assign new_n245_ = new_n232_ & pi018;
  assign new_n246_ = new_n232_ & pi019;
  assign new_n247_ = new_n232_ & pi020;
  assign new_n248_ = new_n232_ & pi021;
  assign new_n249_ = new_n232_ & pi022;
  assign new_n250_ = new_n232_ & pi023;
  assign new_n251_ = new_n232_ & pi024;
  assign new_n252_ = new_n232_ & pi025;
  assign new_n253_ = new_n232_ & pi026;
  assign new_n254_ = new_n232_ & pi027;
  assign new_n255_ = new_n232_ & pi028;
  assign new_n256_ = new_n232_ & pi029;
  assign new_n257_ = new_n232_ & pi030;
  assign new_n258_ = new_n232_ & pi031;
  assign new_n259_ = new_n232_ & pi032;
  assign new_n260_ = new_n232_ & pi033;
  assign new_n261_ = new_n232_ & pi034;
  assign new_n262_ = new_n232_ & pi035;
  assign new_n263_ = new_n232_ & pi036;
  assign new_n264_ = new_n232_ & pi037;
  assign new_n265_ = new_n232_ & pi038;
  assign new_n266_ = new_n232_ & pi039;
  assign new_n267_ = ~new_n232_;
  assign new_n268_ = new_n267_ & pi017 & new_n233_;
  assign new_n269_ = new_n324_ | new_n236_ | new_n268_ | new_n356_ | new_n388_;
  assign new_n270_ = new_n267_ & pi018 & new_n233_;
  assign new_n271_ = new_n325_ | new_n237_ | new_n270_ | new_n357_ | new_n388_;
  assign new_n272_ = new_n267_ & pi019 & new_n233_;
  assign new_n273_ = new_n326_ | new_n238_ | new_n272_ | new_n358_ | new_n388_;
  assign new_n274_ = new_n267_ & pi020 & new_n233_;
  assign new_n275_ = new_n327_ | new_n239_ | new_n274_ | new_n359_ | new_n388_;
  assign new_n276_ = new_n267_ & pi021 & new_n233_;
  assign new_n277_ = new_n328_ | new_n240_ | new_n276_ | new_n360_ | new_n388_;
  assign new_n278_ = new_n267_ & pi022 & new_n233_;
  assign new_n279_ = new_n329_ | new_n241_ | new_n278_ | new_n361_ | new_n388_;
  assign new_n280_ = new_n267_ & pi023 & new_n233_;
  assign new_n281_ = new_n330_ | new_n242_ | new_n280_ | new_n362_ | new_n388_;
  assign new_n282_ = new_n267_ & pi024 & new_n233_;
  assign new_n283_ = new_n331_ | new_n243_ | new_n282_ | new_n363_ | new_n388_;
  assign new_n284_ = new_n267_ & pi025 & new_n233_;
  assign new_n285_ = new_n332_ | new_n244_ | new_n284_ | new_n364_ | new_n388_;
  assign new_n286_ = new_n267_ & pi026 & new_n233_;
  assign new_n287_ = new_n333_ | new_n245_ | new_n286_ | new_n365_ | new_n388_;
  assign new_n288_ = new_n267_ & pi027 & new_n233_;
  assign new_n289_ = new_n334_ | new_n246_ | new_n288_ | new_n366_ | new_n388_;
  assign new_n290_ = new_n267_ & pi028 & new_n233_;
  assign new_n291_ = new_n335_ | new_n247_ | new_n290_ | new_n367_ | new_n388_;
  assign new_n292_ = new_n267_ & pi029 & new_n233_;
  assign new_n293_ = new_n336_ | new_n248_ | new_n292_ | new_n368_ | new_n388_;
  assign new_n294_ = new_n267_ & pi030 & new_n233_;
  assign new_n295_ = new_n337_ | new_n249_ | new_n294_ | new_n369_ | new_n388_;
  assign new_n296_ = new_n267_ & pi031 & new_n233_;
  assign new_n297_ = new_n338_ | new_n250_ | new_n296_ | new_n370_ | new_n388_;
  assign new_n298_ = new_n267_ & pi032 & new_n233_;
  assign new_n299_ = new_n339_ | new_n251_ | new_n298_ | new_n371_ | new_n388_;
  assign new_n300_ = new_n267_ & pi033 & new_n233_;
  assign new_n301_ = new_n340_ | new_n252_ | new_n300_ | new_n372_ | new_n388_;
  assign new_n302_ = new_n267_ & pi034 & new_n233_;
  assign new_n303_ = new_n341_ | new_n253_ | new_n302_ | new_n373_ | new_n388_;
  assign new_n304_ = new_n267_ & pi035 & new_n233_;
  assign new_n305_ = new_n342_ | new_n254_ | new_n304_ | new_n374_ | new_n388_;
  assign new_n306_ = new_n267_ & pi036 & new_n233_;
  assign new_n307_ = new_n343_ | new_n255_ | new_n306_ | new_n375_ | new_n388_;
  assign new_n308_ = new_n267_ & pi037 & new_n233_;
  assign new_n309_ = new_n344_ | new_n256_ | new_n308_ | new_n376_ | new_n388_;
  assign new_n310_ = new_n267_ & pi038 & new_n233_;
  assign new_n311_ = new_n345_ | new_n257_ | new_n310_ | new_n377_ | new_n388_;
  assign new_n312_ = new_n267_ & pi039 & new_n233_;
  assign new_n313_ = new_n346_ | new_n258_ | new_n312_ | new_n378_ | new_n388_;
  assign new_n314_ = new_n267_ & pi040 & new_n233_;
  assign new_n315_ = new_n347_ | new_n259_ | new_n314_ | new_n379_ | new_n388_;
  assign new_n316_ = new_n260_ | new_n388_ | new_n348_ | new_n380_;
  assign new_n317_ = new_n261_ | new_n388_ | new_n349_ | new_n381_;
  assign new_n318_ = new_n262_ | new_n388_ | new_n350_ | new_n382_;
  assign new_n319_ = new_n263_ | new_n388_ | new_n351_ | new_n383_;
  assign new_n320_ = new_n264_ | new_n388_ | new_n352_ | new_n384_;
  assign new_n321_ = new_n265_ | new_n388_ | new_n353_ | new_n385_;
  assign new_n322_ = new_n266_ | new_n388_ | new_n354_ | new_n386_;
  assign new_n323_ = ~new_n233_;
  assign new_n324_ = new_n234_ & new_n267_ & pi020 & new_n323_;
  assign new_n325_ = new_n234_ & new_n267_ & pi021 & new_n323_;
  assign new_n326_ = new_n234_ & new_n267_ & pi022 & new_n323_;
  assign new_n327_ = new_n234_ & new_n267_ & pi023 & new_n323_;
  assign new_n328_ = new_n234_ & new_n267_ & pi024 & new_n323_;
  assign new_n329_ = new_n234_ & new_n267_ & pi025 & new_n323_;
  assign new_n330_ = new_n234_ & new_n267_ & pi026 & new_n323_;
  assign new_n331_ = new_n234_ & new_n267_ & pi027 & new_n323_;
  assign new_n332_ = new_n234_ & new_n267_ & pi028 & new_n323_;
  assign new_n333_ = new_n234_ & new_n267_ & pi029 & new_n323_;
  assign new_n334_ = new_n234_ & new_n267_ & pi030 & new_n323_;
  assign new_n335_ = new_n234_ & new_n267_ & pi031 & new_n323_;
  assign new_n336_ = new_n234_ & new_n267_ & pi032 & new_n323_;
  assign new_n337_ = new_n234_ & new_n267_ & pi033 & new_n323_;
  assign new_n338_ = new_n234_ & new_n267_ & pi034 & new_n323_;
  assign new_n339_ = new_n234_ & new_n267_ & pi035 & new_n323_;
  assign new_n340_ = new_n234_ & new_n267_ & pi036 & new_n323_;
  assign new_n341_ = new_n234_ & new_n267_ & pi037 & new_n323_;
  assign new_n342_ = new_n234_ & new_n267_ & pi038 & new_n323_;
  assign new_n343_ = new_n234_ & new_n267_ & pi039 & new_n323_;
  assign new_n344_ = new_n234_ & new_n267_ & pi041 & new_n323_;
  assign new_n345_ = new_n234_ & new_n267_ & pi042 & new_n323_;
  assign new_n346_ = new_n234_ & new_n267_ & pi043 & new_n323_;
  assign new_n347_ = new_n234_ & new_n267_ & pi044 & new_n323_;
  assign new_n348_ = new_n234_ & new_n267_ & pi045 & new_n323_;
  assign new_n349_ = new_n234_ & new_n267_ & pi046 & new_n323_;
  assign new_n350_ = new_n234_ & new_n267_ & pi047 & new_n323_;
  assign new_n351_ = new_n234_ & new_n267_ & pi048 & new_n323_;
  assign new_n352_ = new_n234_ & new_n267_ & pi049 & new_n323_;
  assign new_n353_ = new_n234_ & new_n267_ & pi050 & new_n323_;
  assign new_n354_ = new_n234_ & new_n267_ & pi051 & new_n323_;
  assign new_n355_ = ~new_n234_;
  assign new_n356_ = new_n235_ & new_n323_ & new_n267_ & pi024 & new_n355_;
  assign new_n357_ = new_n235_ & new_n323_ & new_n267_ & pi025 & new_n355_;
  assign new_n358_ = new_n235_ & new_n323_ & new_n267_ & pi026 & new_n355_;
  assign new_n359_ = new_n235_ & new_n323_ & new_n267_ & pi027 & new_n355_;
  assign new_n360_ = new_n235_ & new_n323_ & new_n267_ & pi028 & new_n355_;
  assign new_n361_ = new_n235_ & new_n323_ & new_n267_ & pi029 & new_n355_;
  assign new_n362_ = new_n235_ & new_n323_ & new_n267_ & pi030 & new_n355_;
  assign new_n363_ = new_n235_ & new_n323_ & new_n267_ & pi031 & new_n355_;
  assign new_n364_ = new_n235_ & new_n323_ & new_n267_ & pi032 & new_n355_;
  assign new_n365_ = new_n235_ & new_n323_ & new_n267_ & pi033 & new_n355_;
  assign new_n366_ = new_n235_ & new_n323_ & new_n267_ & pi034 & new_n355_;
  assign new_n367_ = new_n235_ & new_n323_ & new_n267_ & pi035 & new_n355_;
  assign new_n368_ = new_n235_ & new_n323_ & new_n267_ & pi036 & new_n355_;
  assign new_n369_ = new_n235_ & new_n323_ & new_n267_ & pi037 & new_n355_;
  assign new_n370_ = new_n235_ & new_n323_ & new_n267_ & pi038 & new_n355_;
  assign new_n371_ = new_n235_ & new_n323_ & new_n267_ & pi039 & new_n355_;
  assign new_n372_ = new_n235_ & new_n323_ & new_n267_ & pi052 & new_n355_;
  assign new_n373_ = new_n235_ & new_n323_ & new_n267_ & pi053 & new_n355_;
  assign new_n374_ = new_n235_ & new_n323_ & new_n267_ & pi054 & new_n355_;
  assign new_n375_ = new_n235_ & new_n323_ & new_n267_ & pi055 & new_n355_;
  assign new_n376_ = new_n235_ & new_n323_ & new_n267_ & pi056 & new_n355_;
  assign new_n377_ = new_n235_ & new_n323_ & new_n267_ & pi057 & new_n355_;
  assign new_n378_ = new_n235_ & new_n323_ & new_n267_ & pi058 & new_n355_;
  assign new_n379_ = new_n235_ & new_n323_ & new_n267_ & pi059 & new_n355_;
  assign new_n380_ = new_n235_ & new_n323_ & new_n267_ & pi060 & new_n355_;
  assign new_n381_ = new_n235_ & new_n323_ & new_n267_ & pi061 & new_n355_;
  assign new_n382_ = new_n235_ & new_n323_ & new_n267_ & pi062 & new_n355_;
  assign new_n383_ = new_n235_ & new_n323_ & new_n267_ & pi063 & new_n355_;
  assign new_n384_ = new_n235_ & new_n323_ & new_n267_ & pi064 & new_n355_;
  assign new_n385_ = new_n235_ & new_n323_ & new_n267_ & pi065 & new_n355_;
  assign new_n386_ = new_n235_ & new_n323_ & new_n267_ & pi066 & new_n355_;
  assign new_n387_ = ~new_n235_;
  assign new_n388_ = new_n355_ & new_n267_ & new_n387_ & new_n323_;
  assign new_n389_ = new_n232_ & pi067;
  assign new_n390_ = new_n232_ & pi068;
  assign new_n391_ = new_n232_ & pi069;
  assign new_n392_ = new_n232_ & pi070;
  assign new_n393_ = new_n232_ & pi071;
  assign new_n394_ = new_n232_ & pi072;
  assign new_n395_ = new_n232_ & pi073;
  assign new_n396_ = new_n232_ & pi074;
  assign new_n397_ = new_n232_ & pi075;
  assign new_n398_ = new_n232_ & pi076;
  assign new_n399_ = new_n232_ & pi077;
  assign new_n400_ = new_n232_ & pi078;
  assign new_n401_ = new_n232_ & pi079;
  assign new_n402_ = new_n232_ & pi080;
  assign new_n403_ = new_n232_ & pi081;
  assign new_n404_ = new_n232_ & pi082;
  assign new_n405_ = new_n232_ & pi083;
  assign new_n406_ = new_n232_ & pi084;
  assign new_n407_ = new_n232_ & pi085;
  assign new_n408_ = new_n232_ & pi086;
  assign new_n409_ = new_n232_ & pi041;
  assign new_n410_ = new_n232_ & pi042;
  assign new_n411_ = new_n232_ & pi043;
  assign new_n412_ = new_n232_ & pi044;
  assign new_n413_ = new_n232_ & pi045;
  assign new_n414_ = new_n232_ & pi046;
  assign new_n415_ = new_n232_ & pi047;
  assign new_n416_ = new_n232_ & pi048;
  assign new_n417_ = new_n232_ & pi049;
  assign new_n418_ = new_n232_ & pi050;
  assign new_n419_ = new_n232_ & pi051;
  assign new_n420_ = new_n232_ & pi087;
  assign new_n421_ = ~new_n232_;
  assign new_n422_ = new_n421_ & pi075 & new_n233_;
  assign new_n423_ = new_n487_ | new_n389_ | new_n422_ | new_n520_ | new_n553_;
  assign new_n424_ = new_n421_ & pi076 & new_n233_;
  assign new_n425_ = new_n488_ | new_n390_ | new_n424_ | new_n521_ | new_n553_;
  assign new_n426_ = new_n421_ & pi077 & new_n233_;
  assign new_n427_ = new_n489_ | new_n391_ | new_n426_ | new_n522_ | new_n553_;
  assign new_n428_ = new_n421_ & pi078 & new_n233_;
  assign new_n429_ = new_n490_ | new_n392_ | new_n428_ | new_n523_ | new_n553_;
  assign new_n430_ = new_n421_ & pi079 & new_n233_;
  assign new_n431_ = new_n491_ | new_n393_ | new_n430_ | new_n524_ | new_n553_;
  assign new_n432_ = new_n421_ & pi080 & new_n233_;
  assign new_n433_ = new_n492_ | new_n394_ | new_n432_ | new_n525_ | new_n553_;
  assign new_n434_ = new_n421_ & pi081 & new_n233_;
  assign new_n435_ = new_n493_ | new_n395_ | new_n434_ | new_n526_ | new_n553_;
  assign new_n436_ = new_n421_ & pi082 & new_n233_;
  assign new_n437_ = new_n494_ | new_n396_ | new_n436_ | new_n527_ | new_n553_;
  assign new_n438_ = new_n421_ & pi083 & new_n233_;
  assign new_n439_ = new_n495_ | new_n397_ | new_n438_ | new_n528_ | new_n553_;
  assign new_n440_ = new_n421_ & pi084 & new_n233_;
  assign new_n441_ = new_n496_ | new_n398_ | new_n440_ | new_n529_ | new_n553_;
  assign new_n442_ = new_n421_ & pi085 & new_n233_;
  assign new_n443_ = new_n497_ | new_n399_ | new_n442_ | new_n530_ | new_n553_;
  assign new_n444_ = new_n421_ & pi086 & new_n233_;
  assign new_n445_ = new_n498_ | new_n400_ | new_n444_ | new_n531_ | new_n553_;
  assign new_n446_ = new_n421_ & pi041 & new_n233_;
  assign new_n447_ = new_n499_ | new_n401_ | new_n446_ | new_n532_ | new_n553_;
  assign new_n448_ = new_n421_ & pi042 & new_n233_;
  assign new_n449_ = new_n500_ | new_n402_ | new_n448_ | new_n533_ | new_n553_;
  assign new_n450_ = new_n421_ & pi043 & new_n233_;
  assign new_n451_ = new_n501_ | new_n403_ | new_n450_ | new_n534_ | new_n553_;
  assign new_n452_ = new_n421_ & pi044 & new_n233_;
  assign new_n453_ = new_n502_ | new_n404_ | new_n452_ | new_n535_ | new_n553_;
  assign new_n454_ = new_n421_ & pi045 & new_n233_;
  assign new_n455_ = new_n503_ | new_n405_ | new_n454_ | new_n536_ | new_n553_;
  assign new_n456_ = new_n421_ & pi046 & new_n233_;
  assign new_n457_ = new_n504_ | new_n406_ | new_n456_ | new_n537_ | new_n553_;
  assign new_n458_ = new_n421_ & pi047 & new_n233_;
  assign new_n459_ = new_n505_ | new_n407_ | new_n458_ | new_n538_ | new_n553_;
  assign new_n460_ = new_n421_ & pi048 & new_n233_;
  assign new_n461_ = new_n506_ | new_n408_ | new_n460_ | new_n539_ | new_n553_;
  assign new_n462_ = new_n421_ & pi049 & new_n233_;
  assign new_n463_ = new_n507_ | new_n409_ | new_n462_ | new_n540_ | new_n553_;
  assign new_n464_ = new_n421_ & pi050 & new_n233_;
  assign new_n465_ = new_n508_ | new_n410_ | new_n464_ | new_n541_ | new_n553_;
  assign new_n466_ = new_n421_ & pi051 & new_n233_;
  assign new_n467_ = new_n509_ | new_n411_ | new_n466_ | new_n542_ | new_n553_;
  assign new_n468_ = new_n421_ & pi087 & new_n233_;
  assign new_n469_ = new_n510_ | new_n412_ | new_n468_ | new_n543_ | new_n553_;
  assign new_n470_ = new_n421_ & pi009 & new_n233_;
  assign new_n471_ = new_n511_ | new_n413_ | new_n470_ | new_n544_ | new_n553_;
  assign new_n472_ = new_n421_ & pi010 & new_n233_;
  assign new_n473_ = new_n512_ | new_n414_ | new_n472_ | new_n545_ | new_n553_;
  assign new_n474_ = new_n421_ & pi011 & new_n233_;
  assign new_n475_ = new_n513_ | new_n415_ | new_n474_ | new_n546_ | new_n553_;
  assign new_n476_ = new_n421_ & pi012 & new_n233_;
  assign new_n477_ = new_n514_ | new_n416_ | new_n476_ | new_n547_ | new_n553_;
  assign new_n478_ = new_n421_ & pi013 & new_n233_;
  assign new_n479_ = new_n515_ | new_n417_ | new_n478_ | new_n548_ | new_n553_;
  assign new_n480_ = new_n421_ & pi014 & new_n233_;
  assign new_n481_ = new_n516_ | new_n418_ | new_n480_ | new_n549_ | new_n553_;
  assign new_n482_ = new_n421_ & pi015 & new_n233_;
  assign new_n483_ = new_n517_ | new_n419_ | new_n482_ | new_n550_ | new_n553_;
  assign new_n484_ = new_n421_ & pi016 & new_n233_;
  assign new_n485_ = new_n518_ | new_n420_ | new_n484_ | new_n551_ | new_n553_;
  assign new_n486_ = ~new_n233_;
  assign new_n487_ = new_n234_ & new_n421_ & pi078 & new_n486_;
  assign new_n488_ = new_n234_ & new_n421_ & pi079 & new_n486_;
  assign new_n489_ = new_n234_ & new_n421_ & pi080 & new_n486_;
  assign new_n490_ = new_n234_ & new_n421_ & pi081 & new_n486_;
  assign new_n491_ = new_n234_ & new_n421_ & pi082 & new_n486_;
  assign new_n492_ = new_n234_ & new_n421_ & pi083 & new_n486_;
  assign new_n493_ = new_n234_ & new_n421_ & pi084 & new_n486_;
  assign new_n494_ = new_n234_ & new_n421_ & pi085 & new_n486_;
  assign new_n495_ = new_n234_ & new_n421_ & pi086 & new_n486_;
  assign new_n496_ = new_n234_ & new_n421_ & pi041 & new_n486_;
  assign new_n497_ = new_n234_ & new_n421_ & pi042 & new_n486_;
  assign new_n498_ = new_n234_ & new_n421_ & pi043 & new_n486_;
  assign new_n499_ = new_n234_ & new_n421_ & pi044 & new_n486_;
  assign new_n500_ = new_n234_ & new_n421_ & pi045 & new_n486_;
  assign new_n501_ = new_n234_ & new_n421_ & pi046 & new_n486_;
  assign new_n502_ = new_n234_ & new_n421_ & pi047 & new_n486_;
  assign new_n503_ = new_n234_ & new_n421_ & pi048 & new_n486_;
  assign new_n504_ = new_n234_ & new_n421_ & pi049 & new_n486_;
  assign new_n505_ = new_n234_ & new_n421_ & pi050 & new_n486_;
  assign new_n506_ = new_n234_ & new_n421_ & pi051 & new_n486_;
  assign new_n507_ = new_n234_ & new_n421_ & pi087 & new_n486_;
  assign new_n508_ = new_n234_ & new_n421_ & pi009 & new_n486_;
  assign new_n509_ = new_n234_ & new_n421_ & pi010 & new_n486_;
  assign new_n510_ = new_n234_ & new_n421_ & pi011 & new_n486_;
  assign new_n511_ = new_n234_ & new_n421_ & pi012 & new_n486_;
  assign new_n512_ = new_n234_ & new_n421_ & pi013 & new_n486_;
  assign new_n513_ = new_n234_ & new_n421_ & pi014 & new_n486_;
  assign new_n514_ = new_n234_ & new_n421_ & pi015 & new_n486_;
  assign new_n515_ = new_n234_ & new_n421_ & pi016 & new_n486_;
  assign new_n516_ = new_n234_ & new_n421_ & pi017 & new_n486_;
  assign new_n517_ = new_n234_ & new_n421_ & pi018 & new_n486_;
  assign new_n518_ = new_n234_ & new_n421_ & pi019 & new_n486_;
  assign new_n519_ = ~new_n234_;
  assign new_n520_ = new_n235_ & new_n486_ & new_n421_ & pi082 & new_n519_;
  assign new_n521_ = new_n235_ & new_n486_ & new_n421_ & pi083 & new_n519_;
  assign new_n522_ = new_n235_ & new_n486_ & new_n421_ & pi084 & new_n519_;
  assign new_n523_ = new_n235_ & new_n486_ & new_n421_ & pi085 & new_n519_;
  assign new_n524_ = new_n235_ & new_n486_ & new_n421_ & pi086 & new_n519_;
  assign new_n525_ = new_n235_ & new_n486_ & new_n421_ & pi041 & new_n519_;
  assign new_n526_ = new_n235_ & new_n486_ & new_n421_ & pi042 & new_n519_;
  assign new_n527_ = new_n235_ & new_n486_ & new_n421_ & pi043 & new_n519_;
  assign new_n528_ = new_n235_ & new_n486_ & new_n421_ & pi044 & new_n519_;
  assign new_n529_ = new_n235_ & new_n486_ & new_n421_ & pi045 & new_n519_;
  assign new_n530_ = new_n235_ & new_n486_ & new_n421_ & pi046 & new_n519_;
  assign new_n531_ = new_n235_ & new_n486_ & new_n421_ & pi047 & new_n519_;
  assign new_n532_ = new_n235_ & new_n486_ & new_n421_ & pi048 & new_n519_;
  assign new_n533_ = new_n235_ & new_n486_ & new_n421_ & pi049 & new_n519_;
  assign new_n534_ = new_n235_ & new_n486_ & new_n421_ & pi050 & new_n519_;
  assign new_n535_ = new_n235_ & new_n486_ & new_n421_ & pi051 & new_n519_;
  assign new_n536_ = new_n235_ & new_n486_ & new_n421_ & pi087 & new_n519_;
  assign new_n537_ = new_n235_ & new_n486_ & new_n421_ & pi009 & new_n519_;
  assign new_n538_ = new_n235_ & new_n486_ & new_n421_ & pi010 & new_n519_;
  assign new_n539_ = new_n235_ & new_n486_ & new_n421_ & pi011 & new_n519_;
  assign new_n540_ = new_n235_ & new_n486_ & new_n421_ & pi012 & new_n519_;
  assign new_n541_ = new_n235_ & new_n486_ & new_n421_ & pi013 & new_n519_;
  assign new_n542_ = new_n235_ & new_n486_ & new_n421_ & pi014 & new_n519_;
  assign new_n543_ = new_n235_ & new_n486_ & new_n421_ & pi015 & new_n519_;
  assign new_n544_ = new_n235_ & new_n486_ & new_n421_ & pi016 & new_n519_;
  assign new_n545_ = new_n235_ & new_n486_ & new_n421_ & pi017 & new_n519_;
  assign new_n546_ = new_n235_ & new_n486_ & new_n421_ & pi018 & new_n519_;
  assign new_n547_ = new_n235_ & new_n486_ & new_n421_ & pi019 & new_n519_;
  assign new_n548_ = new_n235_ & new_n486_ & new_n421_ & pi020 & new_n519_;
  assign new_n549_ = new_n235_ & new_n486_ & new_n421_ & pi021 & new_n519_;
  assign new_n550_ = new_n235_ & new_n486_ & new_n421_ & pi022 & new_n519_;
  assign new_n551_ = new_n235_ & new_n486_ & new_n421_ & pi023 & new_n519_;
  assign new_n552_ = ~new_n235_;
  assign new_n553_ = new_n519_ & new_n421_ & new_n552_ & new_n486_;
  assign new_n554_ = new_n1190_ & pi088;
  assign new_n555_ = ~new_n1190_;
  assign new_n556_ = new_n555_ & pi088 & new_n1194_;
  assign po00 = new_n559_ | new_n554_ | new_n556_ | new_n565_ | new_n561_ | new_n563_;
  assign new_n558_ = ~new_n1194_;
  assign new_n559_ = new_n1198_ & new_n555_ & pi089 & new_n558_;
  assign new_n560_ = ~new_n1198_;
  assign new_n561_ = new_n1200_ & new_n558_ & new_n555_ & pi090 & new_n560_;
  assign new_n562_ = ~new_n1200_;
  assign new_n563_ = pi005 & new_n560_ & new_n555_ & new_n558_ & pi087 & new_n562_;
  assign new_n564_ = ~pi005;
  assign new_n565_ = new_n562_ & new_n558_ & new_n555_ & new_n564_ & new_n560_;
  assign new_n566_ = new_n1204_ & new_n321_;
  assign new_n567_ = new_n1204_ & new_n322_;
  assign new_n568_ = ~new_n1204_;
  assign new_n569_ = new_n568_ & new_n321_ & new_n1207_;
  assign po01 = new_n574_ | new_n566_ | new_n569_ | new_n582_ | new_n585_ | new_n579_;
  assign new_n571_ = new_n568_ & new_n322_ & new_n1207_;
  assign po02 = new_n567_ | new_n571_ | new_n575_ | new_n577_ | new_n586_ | new_n580_ | new_n583_;
  assign new_n573_ = ~new_n1207_;
  assign new_n574_ = pi005 & new_n568_ & new_n321_ & new_n573_;
  assign new_n575_ = pi005 & new_n568_ & new_n322_ & new_n573_;
  assign new_n576_ = ~pi005;
  assign new_n577_ = new_n1210_ & new_n573_ & new_n568_ & pi091 & new_n576_;
  assign new_n578_ = ~new_n1210_;
  assign new_n579_ = new_n1215_ & new_n576_ & new_n568_ & new_n573_ & pi092 & new_n578_;
  assign new_n580_ = new_n1215_ & new_n576_ & new_n568_ & new_n573_ & pi093 & new_n578_;
  assign new_n581_ = ~new_n1215_;
  assign new_n582_ = new_n1220_ & new_n578_ & new_n573_ & new_n568_ & new_n576_ & pi092 & new_n581_;
  assign new_n583_ = new_n1220_ & new_n578_ & new_n573_ & new_n568_ & new_n576_ & pi093 & new_n581_;
  assign new_n584_ = ~new_n1220_;
  assign new_n585_ = new_n1221_ & pi095 & new_n581_ & new_n576_ & new_n568_ & new_n573_ & new_n578_ & pi094 & new_n584_;
  assign new_n586_ = new_n1221_ & pi095 & new_n581_ & new_n576_ & new_n568_ & new_n573_ & new_n578_ & pi096 & new_n584_;
  assign new_n587_ = new_n1225_ & new_n315_;
  assign new_n588_ = new_n1225_ & new_n316_;
  assign new_n589_ = new_n1225_ & new_n317_;
  assign new_n590_ = new_n1225_ & new_n318_;
  assign new_n591_ = new_n1225_ & new_n319_;
  assign new_n592_ = new_n1225_ & new_n320_;
  assign new_n593_ = ~new_n1225_;
  assign new_n594_ = new_n593_ & new_n315_ & new_n1227_;
  assign po03 = new_n587_ | new_n594_ | new_n607_ | new_n614_;
  assign new_n596_ = new_n593_ & new_n316_ & new_n1227_;
  assign po04 = new_n588_ | new_n596_ | new_n608_ | new_n615_;
  assign new_n598_ = new_n593_ & new_n317_ & new_n1227_;
  assign po05 = new_n589_ | new_n598_ | new_n609_ | new_n616_;
  assign new_n600_ = new_n593_ & new_n318_ & new_n1227_;
  assign po06 = new_n590_ | new_n600_ | new_n610_ | new_n617_;
  assign new_n602_ = new_n593_ & new_n319_ & new_n1227_;
  assign po07 = new_n591_ | new_n602_ | new_n611_ | new_n618_;
  assign new_n604_ = new_n593_ & new_n320_ & new_n1227_;
  assign po08 = new_n592_ | new_n604_ | new_n612_ | new_n619_;
  assign new_n606_ = ~new_n1227_;
  assign new_n607_ = pi005 & new_n593_ & new_n315_ & new_n606_;
  assign new_n608_ = pi005 & new_n593_ & new_n316_ & new_n606_;
  assign new_n609_ = pi005 & new_n593_ & new_n317_ & new_n606_;
  assign new_n610_ = pi005 & new_n593_ & new_n318_ & new_n606_;
  assign new_n611_ = pi005 & new_n593_ & new_n319_ & new_n606_;
  assign new_n612_ = pi005 & new_n593_ & new_n320_ & new_n606_;
  assign new_n613_ = ~pi005;
  assign new_n614_ = new_n1228_ & pi095 & new_n606_ & new_n593_ & pi097 & new_n613_;
  assign new_n615_ = new_n1228_ & pi095 & new_n606_ & new_n593_ & pi098 & new_n613_;
  assign new_n616_ = new_n1228_ & pi095 & new_n606_ & new_n593_ & pi099 & new_n613_;
  assign new_n617_ = new_n1228_ & pi095 & new_n606_ & new_n593_ & pi100 & new_n613_;
  assign new_n618_ = new_n1228_ & pi095 & new_n606_ & new_n593_ & pi101 & new_n613_;
  assign new_n619_ = new_n1228_ & pi095 & new_n606_ & new_n593_ & pi102 & new_n613_;
  assign new_n620_ = new_n1231_ & new_n313_;
  assign new_n621_ = ~new_n1231_;
  assign new_n622_ = new_n621_ & new_n313_ & new_n1233_;
  assign po09 = new_n620_ | new_n622_ | new_n625_ | new_n627_;
  assign new_n624_ = ~new_n1233_;
  assign new_n625_ = pi005 & new_n621_ & new_n313_ & new_n624_;
  assign new_n626_ = ~pi005;
  assign new_n627_ = new_n1234_ & pi095 & new_n624_ & new_n621_ & pi103 & new_n626_;
  assign new_n628_ = new_n1238_ & new_n309_;
  assign new_n629_ = new_n1238_ & new_n311_;
  assign new_n630_ = ~new_n1238_;
  assign new_n631_ = new_n630_ & new_n309_ & new_n1240_;
  assign po10 = new_n628_ | new_n631_ | new_n636_ | new_n639_;
  assign new_n633_ = new_n630_ & new_n311_ & new_n1240_;
  assign po11 = new_n629_ | new_n633_ | new_n637_ | new_n640_;
  assign new_n635_ = ~new_n1240_;
  assign new_n636_ = pi005 & new_n630_ & new_n309_ & new_n635_;
  assign new_n637_ = pi005 & new_n630_ & new_n311_ & new_n635_;
  assign new_n638_ = ~pi005;
  assign new_n639_ = new_n1241_ & pi095 & new_n635_ & new_n630_ & pi104 & new_n638_;
  assign new_n640_ = new_n1241_ & pi095 & new_n635_ & new_n630_ & pi105 & new_n638_;
  assign new_n641_ = new_n1245_ & new_n307_;
  assign new_n642_ = ~new_n1245_;
  assign new_n643_ = new_n642_ & new_n307_ & new_n1250_;
  assign po12 = new_n641_ | new_n643_ | new_n646_ | new_n648_ | new_n654_ | new_n650_ | new_n652_;
  assign new_n645_ = ~new_n1250_;
  assign new_n646_ = new_n1253_ & new_n642_ & new_n307_ & new_n645_;
  assign new_n647_ = ~new_n1253_;
  assign new_n648_ = new_n1255_ & new_n645_ & new_n642_ & new_n307_ & new_n647_;
  assign new_n649_ = ~new_n1255_;
  assign new_n650_ = pi005 & new_n647_ & new_n642_ & new_n645_ & new_n307_ & new_n649_;
  assign new_n651_ = ~pi005;
  assign new_n652_ = new_n1257_ & new_n649_ & new_n645_ & new_n642_ & new_n647_ & pi106 & new_n651_;
  assign new_n653_ = ~new_n1257_;
  assign new_n654_ = new_n1262_ & pi001 & pi002 & new_n1258_ & new_n1259_ & new_n1261_ & new_n1260_ & new_n651_ & new_n647_ & new_n642_ & new_n645_ & new_n649_ & pi086 & new_n653_;
  assign new_n655_ = new_n1267_ & new_n301_;
  assign new_n656_ = new_n1267_ & new_n303_;
  assign new_n657_ = new_n1267_ & new_n305_;
  assign new_n658_ = ~new_n1267_;
  assign new_n659_ = new_n658_ & new_n301_ & new_n1272_;
  assign po13 = new_n655_ | new_n659_ | new_n666_ | new_n670_ | new_n682_ | new_n674_ | new_n678_;
  assign new_n661_ = new_n658_ & new_n303_ & new_n1272_;
  assign po14 = new_n656_ | new_n661_ | new_n667_ | new_n671_ | new_n683_ | new_n675_ | new_n679_;
  assign new_n663_ = new_n658_ & new_n305_ & new_n1272_;
  assign po15 = new_n657_ | new_n663_ | new_n668_ | new_n672_ | new_n684_ | new_n676_ | new_n680_;
  assign new_n665_ = ~new_n1272_;
  assign new_n666_ = new_n1275_ & new_n658_ & new_n301_ & new_n665_;
  assign new_n667_ = new_n1275_ & new_n658_ & new_n303_ & new_n665_;
  assign new_n668_ = new_n1275_ & new_n658_ & new_n305_ & new_n665_;
  assign new_n669_ = ~new_n1275_;
  assign new_n670_ = new_n1277_ & new_n665_ & new_n658_ & new_n301_ & new_n669_;
  assign new_n671_ = new_n1277_ & new_n665_ & new_n658_ & new_n303_ & new_n669_;
  assign new_n672_ = new_n1277_ & new_n665_ & new_n658_ & new_n305_ & new_n669_;
  assign new_n673_ = ~new_n1277_;
  assign new_n674_ = pi005 & new_n669_ & new_n658_ & new_n665_ & new_n301_ & new_n673_;
  assign new_n675_ = pi005 & new_n669_ & new_n658_ & new_n665_ & new_n303_ & new_n673_;
  assign new_n676_ = pi005 & new_n669_ & new_n658_ & new_n665_ & new_n305_ & new_n673_;
  assign new_n677_ = ~pi005;
  assign new_n678_ = new_n1279_ & new_n673_ & new_n665_ & new_n658_ & new_n669_ & pi107 & new_n677_;
  assign new_n679_ = new_n1279_ & new_n673_ & new_n665_ & new_n658_ & new_n669_ & pi108 & new_n677_;
  assign new_n680_ = new_n1279_ & new_n673_ & new_n665_ & new_n658_ & new_n669_ & pi109 & new_n677_;
  assign new_n681_ = ~new_n1279_;
  assign new_n682_ = new_n1284_ & pi001 & pi002 & new_n1280_ & new_n1281_ & new_n1283_ & new_n1282_ & new_n677_ & new_n669_ & new_n658_ & new_n665_ & new_n673_ & pi083 & new_n681_;
  assign new_n683_ = new_n1284_ & pi001 & pi002 & new_n1280_ & new_n1281_ & new_n1283_ & new_n1282_ & new_n677_ & new_n669_ & new_n658_ & new_n665_ & new_n673_ & pi084 & new_n681_;
  assign new_n684_ = new_n1284_ & pi001 & pi002 & new_n1280_ & new_n1281_ & new_n1283_ & new_n1282_ & new_n677_ & new_n669_ & new_n658_ & new_n665_ & new_n673_ & pi085 & new_n681_;
  assign new_n685_ = new_n1289_ & new_n299_;
  assign new_n686_ = ~new_n1289_;
  assign new_n687_ = new_n686_ & new_n299_ & new_n1294_;
  assign po16 = new_n685_ | new_n687_ | new_n690_ | new_n692_ | new_n694_ | new_n696_ | new_n698_ | new_n700_;
  assign new_n689_ = ~new_n1294_;
  assign new_n690_ = new_n1299_ & new_n686_ & new_n299_ & new_n689_;
  assign new_n691_ = ~new_n1299_;
  assign new_n692_ = new_n1302_ & new_n689_ & new_n686_ & new_n299_ & new_n691_;
  assign new_n693_ = ~new_n1302_;
  assign new_n694_ = new_n1304_ & new_n691_ & new_n686_ & new_n689_ & new_n299_ & new_n693_;
  assign new_n695_ = ~new_n1304_;
  assign new_n696_ = pi005 & new_n693_ & new_n689_ & new_n686_ & new_n691_ & new_n299_ & new_n695_;
  assign new_n697_ = ~pi005;
  assign new_n698_ = new_n1306_ & new_n695_ & new_n691_ & new_n686_ & new_n689_ & new_n693_ & pi110 & new_n697_;
  assign new_n699_ = ~new_n1306_;
  assign new_n700_ = new_n1311_ & pi001 & pi002 & new_n1307_ & new_n1308_ & new_n1310_ & new_n1309_ & new_n697_ & new_n693_ & new_n689_ & new_n686_ & new_n691_ & new_n695_ & pi082 & new_n699_;
  assign new_n701_ = new_n1316_ & new_n269_;
  assign new_n702_ = new_n1316_ & new_n271_;
  assign new_n703_ = new_n1316_ & new_n273_;
  assign new_n704_ = new_n1316_ & new_n275_;
  assign new_n705_ = new_n1316_ & new_n277_;
  assign new_n706_ = new_n1316_ & new_n279_;
  assign new_n707_ = new_n1316_ & new_n281_;
  assign new_n708_ = new_n1316_ & new_n283_;
  assign new_n709_ = new_n1316_ & new_n285_;
  assign new_n710_ = new_n1316_ & new_n287_;
  assign new_n711_ = new_n1316_ & new_n289_;
  assign new_n712_ = new_n1316_ & new_n291_;
  assign new_n713_ = new_n1316_ & new_n293_;
  assign new_n714_ = new_n1316_ & new_n295_;
  assign new_n715_ = new_n1316_ & new_n297_;
  assign new_n716_ = ~new_n1316_;
  assign new_n717_ = new_n716_ & new_n269_ & new_n1321_;
  assign po17 = new_n701_ | new_n717_ | new_n748_ | new_n764_ | new_n812_ | new_n780_ | new_n796_;
  assign new_n719_ = new_n716_ & new_n271_ & new_n1321_;
  assign po18 = new_n702_ | new_n719_ | new_n749_ | new_n765_ | new_n813_ | new_n781_ | new_n797_;
  assign new_n721_ = new_n716_ & new_n273_ & new_n1321_;
  assign po19 = new_n703_ | new_n721_ | new_n750_ | new_n766_ | new_n814_ | new_n782_ | new_n798_;
  assign new_n723_ = new_n716_ & new_n275_ & new_n1321_;
  assign po20 = new_n704_ | new_n723_ | new_n751_ | new_n767_ | new_n815_ | new_n783_ | new_n799_;
  assign new_n725_ = new_n716_ & new_n277_ & new_n1321_;
  assign po21 = new_n705_ | new_n725_ | new_n752_ | new_n768_ | new_n816_ | new_n784_ | new_n800_;
  assign new_n727_ = new_n716_ & new_n279_ & new_n1321_;
  assign po22 = new_n706_ | new_n727_ | new_n753_ | new_n769_ | new_n817_ | new_n785_ | new_n801_;
  assign new_n729_ = new_n716_ & new_n281_ & new_n1321_;
  assign po23 = new_n707_ | new_n729_ | new_n754_ | new_n770_ | new_n818_ | new_n786_ | new_n802_;
  assign new_n731_ = new_n716_ & new_n283_ & new_n1321_;
  assign po24 = new_n708_ | new_n731_ | new_n755_ | new_n771_ | new_n819_ | new_n787_ | new_n803_;
  assign new_n733_ = new_n716_ & new_n285_ & new_n1321_;
  assign po25 = new_n709_ | new_n733_ | new_n756_ | new_n772_ | new_n820_ | new_n788_ | new_n804_;
  assign new_n735_ = new_n716_ & new_n287_ & new_n1321_;
  assign po26 = new_n710_ | new_n735_ | new_n757_ | new_n773_ | new_n821_ | new_n789_ | new_n805_;
  assign new_n737_ = new_n716_ & new_n289_ & new_n1321_;
  assign po27 = new_n711_ | new_n737_ | new_n758_ | new_n774_ | new_n822_ | new_n790_ | new_n806_;
  assign new_n739_ = new_n716_ & new_n291_ & new_n1321_;
  assign po28 = new_n712_ | new_n739_ | new_n759_ | new_n775_ | new_n823_ | new_n791_ | new_n807_;
  assign new_n741_ = new_n716_ & new_n293_ & new_n1321_;
  assign po29 = new_n713_ | new_n741_ | new_n760_ | new_n776_ | new_n824_ | new_n792_ | new_n808_;
  assign new_n743_ = new_n716_ & new_n295_ & new_n1321_;
  assign po30 = new_n714_ | new_n743_ | new_n761_ | new_n777_ | new_n825_ | new_n793_ | new_n809_;
  assign new_n745_ = new_n716_ & new_n297_ & new_n1321_;
  assign po31 = new_n715_ | new_n745_ | new_n762_ | new_n778_ | new_n826_ | new_n794_ | new_n810_;
  assign new_n747_ = ~new_n1321_;
  assign new_n748_ = new_n1324_ & new_n716_ & new_n269_ & new_n747_;
  assign new_n749_ = new_n1324_ & new_n716_ & new_n271_ & new_n747_;
  assign new_n750_ = new_n1324_ & new_n716_ & new_n273_ & new_n747_;
  assign new_n751_ = new_n1324_ & new_n716_ & new_n275_ & new_n747_;
  assign new_n752_ = new_n1324_ & new_n716_ & new_n277_ & new_n747_;
  assign new_n753_ = new_n1324_ & new_n716_ & new_n279_ & new_n747_;
  assign new_n754_ = new_n1324_ & new_n716_ & new_n281_ & new_n747_;
  assign new_n755_ = new_n1324_ & new_n716_ & new_n283_ & new_n747_;
  assign new_n756_ = new_n1324_ & new_n716_ & new_n285_ & new_n747_;
  assign new_n757_ = new_n1324_ & new_n716_ & new_n287_ & new_n747_;
  assign new_n758_ = new_n1324_ & new_n716_ & new_n289_ & new_n747_;
  assign new_n759_ = new_n1324_ & new_n716_ & new_n291_ & new_n747_;
  assign new_n760_ = new_n1324_ & new_n716_ & new_n293_ & new_n747_;
  assign new_n761_ = new_n1324_ & new_n716_ & new_n295_ & new_n747_;
  assign new_n762_ = new_n1324_ & new_n716_ & new_n297_ & new_n747_;
  assign new_n763_ = ~new_n1324_;
  assign new_n764_ = new_n1326_ & new_n747_ & new_n716_ & new_n269_ & new_n763_;
  assign new_n765_ = new_n1326_ & new_n747_ & new_n716_ & new_n271_ & new_n763_;
  assign new_n766_ = new_n1326_ & new_n747_ & new_n716_ & new_n273_ & new_n763_;
  assign new_n767_ = new_n1326_ & new_n747_ & new_n716_ & new_n275_ & new_n763_;
  assign new_n768_ = new_n1326_ & new_n747_ & new_n716_ & new_n277_ & new_n763_;
  assign new_n769_ = new_n1326_ & new_n747_ & new_n716_ & new_n279_ & new_n763_;
  assign new_n770_ = new_n1326_ & new_n747_ & new_n716_ & new_n281_ & new_n763_;
  assign new_n771_ = new_n1326_ & new_n747_ & new_n716_ & new_n283_ & new_n763_;
  assign new_n772_ = new_n1326_ & new_n747_ & new_n716_ & new_n285_ & new_n763_;
  assign new_n773_ = new_n1326_ & new_n747_ & new_n716_ & new_n287_ & new_n763_;
  assign new_n774_ = new_n1326_ & new_n747_ & new_n716_ & new_n289_ & new_n763_;
  assign new_n775_ = new_n1326_ & new_n747_ & new_n716_ & new_n291_ & new_n763_;
  assign new_n776_ = new_n1326_ & new_n747_ & new_n716_ & new_n293_ & new_n763_;
  assign new_n777_ = new_n1326_ & new_n747_ & new_n716_ & new_n295_ & new_n763_;
  assign new_n778_ = new_n1326_ & new_n747_ & new_n716_ & new_n297_ & new_n763_;
  assign new_n779_ = ~new_n1326_;
  assign new_n780_ = pi005 & new_n763_ & new_n716_ & new_n747_ & new_n269_ & new_n779_;
  assign new_n781_ = pi005 & new_n763_ & new_n716_ & new_n747_ & new_n271_ & new_n779_;
  assign new_n782_ = pi005 & new_n763_ & new_n716_ & new_n747_ & new_n273_ & new_n779_;
  assign new_n783_ = pi005 & new_n763_ & new_n716_ & new_n747_ & new_n275_ & new_n779_;
  assign new_n784_ = pi005 & new_n763_ & new_n716_ & new_n747_ & new_n277_ & new_n779_;
  assign new_n785_ = pi005 & new_n763_ & new_n716_ & new_n747_ & new_n279_ & new_n779_;
  assign new_n786_ = pi005 & new_n763_ & new_n716_ & new_n747_ & new_n281_ & new_n779_;
  assign new_n787_ = pi005 & new_n763_ & new_n716_ & new_n747_ & new_n283_ & new_n779_;
  assign new_n788_ = pi005 & new_n763_ & new_n716_ & new_n747_ & new_n285_ & new_n779_;
  assign new_n789_ = pi005 & new_n763_ & new_n716_ & new_n747_ & new_n287_ & new_n779_;
  assign new_n790_ = pi005 & new_n763_ & new_n716_ & new_n747_ & new_n289_ & new_n779_;
  assign new_n791_ = pi005 & new_n763_ & new_n716_ & new_n747_ & new_n291_ & new_n779_;
  assign new_n792_ = pi005 & new_n763_ & new_n716_ & new_n747_ & new_n293_ & new_n779_;
  assign new_n793_ = pi005 & new_n763_ & new_n716_ & new_n747_ & new_n295_ & new_n779_;
  assign new_n794_ = pi005 & new_n763_ & new_n716_ & new_n747_ & new_n297_ & new_n779_;
  assign new_n795_ = ~pi005;
  assign new_n796_ = new_n1328_ & new_n779_ & new_n747_ & new_n716_ & new_n763_ & pi111 & new_n795_;
  assign new_n797_ = new_n1328_ & new_n779_ & new_n747_ & new_n716_ & new_n763_ & pi112 & new_n795_;
  assign new_n798_ = new_n1328_ & new_n779_ & new_n747_ & new_n716_ & new_n763_ & pi113 & new_n795_;
  assign new_n799_ = new_n1328_ & new_n779_ & new_n747_ & new_n716_ & new_n763_ & pi114 & new_n795_;
  assign new_n800_ = new_n1328_ & new_n779_ & new_n747_ & new_n716_ & new_n763_ & pi115 & new_n795_;
  assign new_n801_ = new_n1328_ & new_n779_ & new_n747_ & new_n716_ & new_n763_ & pi116 & new_n795_;
  assign new_n802_ = new_n1328_ & new_n779_ & new_n747_ & new_n716_ & new_n763_ & pi117 & new_n795_;
  assign new_n803_ = new_n1328_ & new_n779_ & new_n747_ & new_n716_ & new_n763_ & pi118 & new_n795_;
  assign new_n804_ = new_n1328_ & new_n779_ & new_n747_ & new_n716_ & new_n763_ & pi119 & new_n795_;
  assign new_n805_ = new_n1328_ & new_n779_ & new_n747_ & new_n716_ & new_n763_ & pi120 & new_n795_;
  assign new_n806_ = new_n1328_ & new_n779_ & new_n747_ & new_n716_ & new_n763_ & pi121 & new_n795_;
  assign new_n807_ = new_n1328_ & new_n779_ & new_n747_ & new_n716_ & new_n763_ & pi122 & new_n795_;
  assign new_n808_ = new_n1328_ & new_n779_ & new_n747_ & new_n716_ & new_n763_ & pi123 & new_n795_;
  assign new_n809_ = new_n1328_ & new_n779_ & new_n747_ & new_n716_ & new_n763_ & pi124 & new_n795_;
  assign new_n810_ = new_n1328_ & new_n779_ & new_n747_ & new_n716_ & new_n763_ & pi125 & new_n795_;
  assign new_n811_ = ~new_n1328_;
  assign new_n812_ = new_n1333_ & pi001 & pi002 & new_n1329_ & new_n1330_ & new_n1332_ & new_n1331_ & new_n795_ & new_n763_ & new_n716_ & new_n747_ & new_n779_ & pi067 & new_n811_;
  assign new_n813_ = new_n1333_ & pi001 & pi002 & new_n1329_ & new_n1330_ & new_n1332_ & new_n1331_ & new_n795_ & new_n763_ & new_n716_ & new_n747_ & new_n779_ & pi068 & new_n811_;
  assign new_n814_ = new_n1333_ & pi001 & pi002 & new_n1329_ & new_n1330_ & new_n1332_ & new_n1331_ & new_n795_ & new_n763_ & new_n716_ & new_n747_ & new_n779_ & pi069 & new_n811_;
  assign new_n815_ = new_n1333_ & pi001 & pi002 & new_n1329_ & new_n1330_ & new_n1332_ & new_n1331_ & new_n795_ & new_n763_ & new_n716_ & new_n747_ & new_n779_ & pi070 & new_n811_;
  assign new_n816_ = new_n1333_ & pi001 & pi002 & new_n1329_ & new_n1330_ & new_n1332_ & new_n1331_ & new_n795_ & new_n763_ & new_n716_ & new_n747_ & new_n779_ & pi071 & new_n811_;
  assign new_n817_ = new_n1333_ & pi001 & pi002 & new_n1329_ & new_n1330_ & new_n1332_ & new_n1331_ & new_n795_ & new_n763_ & new_n716_ & new_n747_ & new_n779_ & pi072 & new_n811_;
  assign new_n818_ = new_n1333_ & pi001 & pi002 & new_n1329_ & new_n1330_ & new_n1332_ & new_n1331_ & new_n795_ & new_n763_ & new_n716_ & new_n747_ & new_n779_ & pi073 & new_n811_;
  assign new_n819_ = new_n1333_ & pi001 & pi002 & new_n1329_ & new_n1330_ & new_n1332_ & new_n1331_ & new_n795_ & new_n763_ & new_n716_ & new_n747_ & new_n779_ & pi074 & new_n811_;
  assign new_n820_ = new_n1333_ & pi001 & pi002 & new_n1329_ & new_n1330_ & new_n1332_ & new_n1331_ & new_n795_ & new_n763_ & new_n716_ & new_n747_ & new_n779_ & pi075 & new_n811_;
  assign new_n821_ = new_n1333_ & pi001 & pi002 & new_n1329_ & new_n1330_ & new_n1332_ & new_n1331_ & new_n795_ & new_n763_ & new_n716_ & new_n747_ & new_n779_ & pi076 & new_n811_;
  assign new_n822_ = new_n1333_ & pi001 & pi002 & new_n1329_ & new_n1330_ & new_n1332_ & new_n1331_ & new_n795_ & new_n763_ & new_n716_ & new_n747_ & new_n779_ & pi077 & new_n811_;
  assign new_n823_ = new_n1333_ & pi001 & pi002 & new_n1329_ & new_n1330_ & new_n1332_ & new_n1331_ & new_n795_ & new_n763_ & new_n716_ & new_n747_ & new_n779_ & pi078 & new_n811_;
  assign new_n824_ = new_n1333_ & pi001 & pi002 & new_n1329_ & new_n1330_ & new_n1332_ & new_n1331_ & new_n795_ & new_n763_ & new_n716_ & new_n747_ & new_n779_ & pi079 & new_n811_;
  assign new_n825_ = new_n1333_ & pi001 & pi002 & new_n1329_ & new_n1330_ & new_n1332_ & new_n1331_ & new_n795_ & new_n763_ & new_n716_ & new_n747_ & new_n779_ & pi080 & new_n811_;
  assign new_n826_ = new_n1333_ & pi001 & pi002 & new_n1329_ & new_n1330_ & new_n1332_ & new_n1331_ & new_n795_ & new_n763_ & new_n716_ & new_n747_ & new_n779_ & pi081 & new_n811_;
  assign new_n827_ = new_n1339_ & new_n423_;
  assign new_n828_ = new_n1339_ & new_n425_;
  assign new_n829_ = new_n1339_ & new_n427_;
  assign new_n830_ = new_n1339_ & new_n429_;
  assign new_n831_ = new_n1339_ & new_n431_;
  assign new_n832_ = new_n1339_ & new_n433_;
  assign new_n833_ = new_n1339_ & new_n435_;
  assign new_n834_ = new_n1339_ & new_n437_;
  assign new_n835_ = new_n1339_ & new_n439_;
  assign new_n836_ = new_n1339_ & new_n441_;
  assign new_n837_ = new_n1339_ & new_n443_;
  assign new_n838_ = new_n1339_ & new_n445_;
  assign new_n839_ = new_n1339_ & new_n447_;
  assign new_n840_ = new_n1339_ & new_n449_;
  assign new_n841_ = new_n1339_ & new_n451_;
  assign new_n842_ = new_n1339_ & new_n453_;
  assign new_n843_ = new_n1339_ & new_n455_;
  assign new_n844_ = new_n1339_ & new_n457_;
  assign new_n845_ = new_n1339_ & new_n459_;
  assign new_n846_ = new_n1339_ & new_n461_;
  assign new_n847_ = new_n1339_ & new_n463_;
  assign new_n848_ = new_n1339_ & new_n465_;
  assign new_n849_ = new_n1339_ & new_n467_;
  assign new_n850_ = new_n1339_ & new_n469_;
  assign new_n851_ = new_n1339_ & new_n471_;
  assign new_n852_ = new_n1339_ & new_n473_;
  assign new_n853_ = new_n1339_ & new_n475_;
  assign new_n854_ = new_n1339_ & new_n477_;
  assign new_n855_ = new_n1339_ & new_n479_;
  assign new_n856_ = new_n1339_ & new_n481_;
  assign new_n857_ = new_n1339_ & new_n483_;
  assign new_n858_ = new_n1339_ & new_n485_;
  assign new_n859_ = ~new_n1339_;
  assign new_n860_ = new_n859_ & new_n423_ & new_n1343_;
  assign po32 = new_n827_ | new_n860_ | new_n925_ | new_n958_ | new_n1057_ | new_n991_ | new_n1024_;
  assign new_n862_ = new_n859_ & new_n425_ & new_n1343_;
  assign po33 = new_n828_ | new_n862_ | new_n926_ | new_n959_ | new_n1058_ | new_n992_ | new_n1025_;
  assign new_n864_ = new_n859_ & new_n427_ & new_n1343_;
  assign po34 = new_n829_ | new_n864_ | new_n927_ | new_n960_ | new_n1059_ | new_n993_ | new_n1026_;
  assign new_n866_ = new_n859_ & new_n429_ & new_n1343_;
  assign po35 = new_n830_ | new_n866_ | new_n928_ | new_n961_ | new_n1060_ | new_n994_ | new_n1027_;
  assign new_n868_ = new_n859_ & new_n431_ & new_n1343_;
  assign po36 = new_n831_ | new_n868_ | new_n929_ | new_n962_ | new_n1061_ | new_n995_ | new_n1028_;
  assign new_n870_ = new_n859_ & new_n433_ & new_n1343_;
  assign po37 = new_n832_ | new_n870_ | new_n930_ | new_n963_ | new_n1062_ | new_n996_ | new_n1029_;
  assign new_n872_ = new_n859_ & new_n435_ & new_n1343_;
  assign po38 = new_n833_ | new_n872_ | new_n931_ | new_n964_ | new_n1063_ | new_n997_ | new_n1030_;
  assign new_n874_ = new_n859_ & new_n437_ & new_n1343_;
  assign po39 = new_n834_ | new_n874_ | new_n932_ | new_n965_ | new_n1064_ | new_n998_ | new_n1031_;
  assign new_n876_ = new_n859_ & new_n439_ & new_n1343_;
  assign po40 = new_n835_ | new_n876_ | new_n933_ | new_n966_ | new_n1065_ | new_n999_ | new_n1032_;
  assign new_n878_ = new_n859_ & new_n441_ & new_n1343_;
  assign po41 = new_n836_ | new_n878_ | new_n934_ | new_n967_ | new_n1066_ | new_n1000_ | new_n1033_;
  assign new_n880_ = new_n859_ & new_n443_ & new_n1343_;
  assign po42 = new_n837_ | new_n880_ | new_n935_ | new_n968_ | new_n1067_ | new_n1001_ | new_n1034_;
  assign new_n882_ = new_n859_ & new_n445_ & new_n1343_;
  assign po43 = new_n838_ | new_n882_ | new_n936_ | new_n969_ | new_n1068_ | new_n1002_ | new_n1035_;
  assign new_n884_ = new_n859_ & new_n447_ & new_n1343_;
  assign po44 = new_n839_ | new_n884_ | new_n937_ | new_n970_ | new_n1069_ | new_n1003_ | new_n1036_;
  assign new_n886_ = new_n859_ & new_n449_ & new_n1343_;
  assign po45 = new_n840_ | new_n886_ | new_n938_ | new_n971_ | new_n1070_ | new_n1004_ | new_n1037_;
  assign new_n888_ = new_n859_ & new_n451_ & new_n1343_;
  assign po46 = new_n841_ | new_n888_ | new_n939_ | new_n972_ | new_n1071_ | new_n1005_ | new_n1038_;
  assign new_n890_ = new_n859_ & new_n453_ & new_n1343_;
  assign po47 = new_n842_ | new_n890_ | new_n940_ | new_n973_ | new_n1072_ | new_n1006_ | new_n1039_;
  assign new_n892_ = new_n859_ & new_n455_ & new_n1343_;
  assign po48 = new_n843_ | new_n892_ | new_n941_ | new_n974_ | new_n1073_ | new_n1007_ | new_n1040_;
  assign new_n894_ = new_n859_ & new_n457_ & new_n1343_;
  assign po49 = new_n844_ | new_n894_ | new_n942_ | new_n975_ | new_n1074_ | new_n1008_ | new_n1041_;
  assign new_n896_ = new_n859_ & new_n459_ & new_n1343_;
  assign po50 = new_n845_ | new_n896_ | new_n943_ | new_n976_ | new_n1075_ | new_n1009_ | new_n1042_;
  assign new_n898_ = new_n859_ & new_n461_ & new_n1343_;
  assign po51 = new_n846_ | new_n898_ | new_n944_ | new_n977_ | new_n1076_ | new_n1010_ | new_n1043_;
  assign new_n900_ = new_n859_ & new_n463_ & new_n1343_;
  assign po52 = new_n847_ | new_n900_ | new_n945_ | new_n978_ | new_n1077_ | new_n1011_ | new_n1044_;
  assign new_n902_ = new_n859_ & new_n465_ & new_n1343_;
  assign po53 = new_n848_ | new_n902_ | new_n946_ | new_n979_ | new_n1078_ | new_n1012_ | new_n1045_;
  assign new_n904_ = new_n859_ & new_n467_ & new_n1343_;
  assign po54 = new_n849_ | new_n904_ | new_n947_ | new_n980_ | new_n1079_ | new_n1013_ | new_n1046_;
  assign new_n906_ = new_n859_ & new_n469_ & new_n1343_;
  assign po55 = new_n850_ | new_n906_ | new_n948_ | new_n981_ | new_n1080_ | new_n1014_ | new_n1047_;
  assign new_n908_ = new_n859_ & new_n471_ & new_n1343_;
  assign po56 = new_n851_ | new_n908_ | new_n949_ | new_n982_ | new_n1081_ | new_n1015_ | new_n1048_;
  assign new_n910_ = new_n859_ & new_n473_ & new_n1343_;
  assign po57 = new_n852_ | new_n910_ | new_n950_ | new_n983_ | new_n1082_ | new_n1016_ | new_n1049_;
  assign new_n912_ = new_n859_ & new_n475_ & new_n1343_;
  assign po58 = new_n853_ | new_n912_ | new_n951_ | new_n984_ | new_n1083_ | new_n1017_ | new_n1050_;
  assign new_n914_ = new_n859_ & new_n477_ & new_n1343_;
  assign po59 = new_n854_ | new_n914_ | new_n952_ | new_n985_ | new_n1084_ | new_n1018_ | new_n1051_;
  assign new_n916_ = new_n859_ & new_n479_ & new_n1343_;
  assign po60 = new_n855_ | new_n916_ | new_n953_ | new_n986_ | new_n1085_ | new_n1019_ | new_n1052_;
  assign new_n918_ = new_n859_ & new_n481_ & new_n1343_;
  assign po61 = new_n856_ | new_n918_ | new_n954_ | new_n987_ | new_n1086_ | new_n1020_ | new_n1053_;
  assign new_n920_ = new_n859_ & new_n483_ & new_n1343_;
  assign po62 = new_n857_ | new_n920_ | new_n955_ | new_n988_ | new_n1087_ | new_n1021_ | new_n1054_;
  assign new_n922_ = new_n859_ & new_n485_ & new_n1343_;
  assign po63 = new_n858_ | new_n922_ | new_n956_ | new_n989_ | new_n1088_ | new_n1022_ | new_n1055_;
  assign new_n924_ = ~new_n1343_;
  assign new_n925_ = new_n1347_ & new_n859_ & new_n423_ & new_n924_;
  assign new_n926_ = new_n1347_ & new_n859_ & new_n425_ & new_n924_;
  assign new_n927_ = new_n1347_ & new_n859_ & new_n427_ & new_n924_;
  assign new_n928_ = new_n1347_ & new_n859_ & new_n429_ & new_n924_;
  assign new_n929_ = new_n1347_ & new_n859_ & new_n431_ & new_n924_;
  assign new_n930_ = new_n1347_ & new_n859_ & new_n433_ & new_n924_;
  assign new_n931_ = new_n1347_ & new_n859_ & new_n435_ & new_n924_;
  assign new_n932_ = new_n1347_ & new_n859_ & new_n437_ & new_n924_;
  assign new_n933_ = new_n1347_ & new_n859_ & new_n439_ & new_n924_;
  assign new_n934_ = new_n1347_ & new_n859_ & new_n441_ & new_n924_;
  assign new_n935_ = new_n1347_ & new_n859_ & new_n443_ & new_n924_;
  assign new_n936_ = new_n1347_ & new_n859_ & new_n445_ & new_n924_;
  assign new_n937_ = new_n1347_ & new_n859_ & new_n447_ & new_n924_;
  assign new_n938_ = new_n1347_ & new_n859_ & new_n449_ & new_n924_;
  assign new_n939_ = new_n1347_ & new_n859_ & new_n451_ & new_n924_;
  assign new_n940_ = new_n1347_ & new_n859_ & new_n453_ & new_n924_;
  assign new_n941_ = new_n1347_ & new_n859_ & new_n455_ & new_n924_;
  assign new_n942_ = new_n1347_ & new_n859_ & new_n457_ & new_n924_;
  assign new_n943_ = new_n1347_ & new_n859_ & new_n459_ & new_n924_;
  assign new_n944_ = new_n1347_ & new_n859_ & new_n461_ & new_n924_;
  assign new_n945_ = new_n1347_ & new_n859_ & new_n463_ & new_n924_;
  assign new_n946_ = new_n1347_ & new_n859_ & new_n465_ & new_n924_;
  assign new_n947_ = new_n1347_ & new_n859_ & new_n467_ & new_n924_;
  assign new_n948_ = new_n1347_ & new_n859_ & new_n469_ & new_n924_;
  assign new_n949_ = new_n1347_ & new_n859_ & new_n471_ & new_n924_;
  assign new_n950_ = new_n1347_ & new_n859_ & new_n473_ & new_n924_;
  assign new_n951_ = new_n1347_ & new_n859_ & new_n475_ & new_n924_;
  assign new_n952_ = new_n1347_ & new_n859_ & new_n477_ & new_n924_;
  assign new_n953_ = new_n1347_ & new_n859_ & new_n479_ & new_n924_;
  assign new_n954_ = new_n1347_ & new_n859_ & new_n481_ & new_n924_;
  assign new_n955_ = new_n1347_ & new_n859_ & new_n483_ & new_n924_;
  assign new_n956_ = new_n1347_ & new_n859_ & new_n485_ & new_n924_;
  assign new_n957_ = ~new_n1347_;
  assign new_n958_ = new_n1351_ & new_n924_ & new_n859_ & new_n423_ & new_n957_;
  assign new_n959_ = new_n1351_ & new_n924_ & new_n859_ & new_n425_ & new_n957_;
  assign new_n960_ = new_n1351_ & new_n924_ & new_n859_ & new_n427_ & new_n957_;
  assign new_n961_ = new_n1351_ & new_n924_ & new_n859_ & new_n429_ & new_n957_;
  assign new_n962_ = new_n1351_ & new_n924_ & new_n859_ & new_n431_ & new_n957_;
  assign new_n963_ = new_n1351_ & new_n924_ & new_n859_ & new_n433_ & new_n957_;
  assign new_n964_ = new_n1351_ & new_n924_ & new_n859_ & new_n435_ & new_n957_;
  assign new_n965_ = new_n1351_ & new_n924_ & new_n859_ & new_n437_ & new_n957_;
  assign new_n966_ = new_n1351_ & new_n924_ & new_n859_ & new_n439_ & new_n957_;
  assign new_n967_ = new_n1351_ & new_n924_ & new_n859_ & new_n441_ & new_n957_;
  assign new_n968_ = new_n1351_ & new_n924_ & new_n859_ & new_n443_ & new_n957_;
  assign new_n969_ = new_n1351_ & new_n924_ & new_n859_ & new_n445_ & new_n957_;
  assign new_n970_ = new_n1351_ & new_n924_ & new_n859_ & new_n447_ & new_n957_;
  assign new_n971_ = new_n1351_ & new_n924_ & new_n859_ & new_n449_ & new_n957_;
  assign new_n972_ = new_n1351_ & new_n924_ & new_n859_ & new_n451_ & new_n957_;
  assign new_n973_ = new_n1351_ & new_n924_ & new_n859_ & new_n453_ & new_n957_;
  assign new_n974_ = new_n1351_ & new_n924_ & new_n859_ & new_n455_ & new_n957_;
  assign new_n975_ = new_n1351_ & new_n924_ & new_n859_ & new_n457_ & new_n957_;
  assign new_n976_ = new_n1351_ & new_n924_ & new_n859_ & new_n459_ & new_n957_;
  assign new_n977_ = new_n1351_ & new_n924_ & new_n859_ & new_n461_ & new_n957_;
  assign new_n978_ = new_n1351_ & new_n924_ & new_n859_ & new_n463_ & new_n957_;
  assign new_n979_ = new_n1351_ & new_n924_ & new_n859_ & new_n465_ & new_n957_;
  assign new_n980_ = new_n1351_ & new_n924_ & new_n859_ & new_n467_ & new_n957_;
  assign new_n981_ = new_n1351_ & new_n924_ & new_n859_ & new_n469_ & new_n957_;
  assign new_n982_ = new_n1351_ & new_n924_ & new_n859_ & new_n471_ & new_n957_;
  assign new_n983_ = new_n1351_ & new_n924_ & new_n859_ & new_n473_ & new_n957_;
  assign new_n984_ = new_n1351_ & new_n924_ & new_n859_ & new_n475_ & new_n957_;
  assign new_n985_ = new_n1351_ & new_n924_ & new_n859_ & new_n477_ & new_n957_;
  assign new_n986_ = new_n1351_ & new_n924_ & new_n859_ & new_n479_ & new_n957_;
  assign new_n987_ = new_n1351_ & new_n924_ & new_n859_ & new_n481_ & new_n957_;
  assign new_n988_ = new_n1351_ & new_n924_ & new_n859_ & new_n483_ & new_n957_;
  assign new_n989_ = new_n1351_ & new_n924_ & new_n859_ & new_n485_ & new_n957_;
  assign new_n990_ = ~new_n1351_;
  assign new_n991_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n423_ & new_n990_;
  assign new_n992_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n425_ & new_n990_;
  assign new_n993_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n427_ & new_n990_;
  assign new_n994_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n429_ & new_n990_;
  assign new_n995_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n431_ & new_n990_;
  assign new_n996_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n433_ & new_n990_;
  assign new_n997_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n435_ & new_n990_;
  assign new_n998_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n437_ & new_n990_;
  assign new_n999_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n439_ & new_n990_;
  assign new_n1000_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n441_ & new_n990_;
  assign new_n1001_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n443_ & new_n990_;
  assign new_n1002_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n445_ & new_n990_;
  assign new_n1003_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n447_ & new_n990_;
  assign new_n1004_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n449_ & new_n990_;
  assign new_n1005_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n451_ & new_n990_;
  assign new_n1006_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n453_ & new_n990_;
  assign new_n1007_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n455_ & new_n990_;
  assign new_n1008_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n457_ & new_n990_;
  assign new_n1009_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n459_ & new_n990_;
  assign new_n1010_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n461_ & new_n990_;
  assign new_n1011_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n463_ & new_n990_;
  assign new_n1012_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n465_ & new_n990_;
  assign new_n1013_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n467_ & new_n990_;
  assign new_n1014_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n469_ & new_n990_;
  assign new_n1015_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n471_ & new_n990_;
  assign new_n1016_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n473_ & new_n990_;
  assign new_n1017_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n475_ & new_n990_;
  assign new_n1018_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n477_ & new_n990_;
  assign new_n1019_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n479_ & new_n990_;
  assign new_n1020_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n481_ & new_n990_;
  assign new_n1021_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n483_ & new_n990_;
  assign new_n1022_ = new_n1354_ & new_n957_ & new_n859_ & new_n924_ & new_n485_ & new_n990_;
  assign new_n1023_ = ~new_n1354_;
  assign new_n1024_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n423_ & new_n1023_;
  assign new_n1025_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n425_ & new_n1023_;
  assign new_n1026_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n427_ & new_n1023_;
  assign new_n1027_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n429_ & new_n1023_;
  assign new_n1028_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n431_ & new_n1023_;
  assign new_n1029_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n433_ & new_n1023_;
  assign new_n1030_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n435_ & new_n1023_;
  assign new_n1031_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n437_ & new_n1023_;
  assign new_n1032_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n439_ & new_n1023_;
  assign new_n1033_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n441_ & new_n1023_;
  assign new_n1034_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n443_ & new_n1023_;
  assign new_n1035_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n445_ & new_n1023_;
  assign new_n1036_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n447_ & new_n1023_;
  assign new_n1037_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n449_ & new_n1023_;
  assign new_n1038_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n451_ & new_n1023_;
  assign new_n1039_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n453_ & new_n1023_;
  assign new_n1040_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n455_ & new_n1023_;
  assign new_n1041_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n457_ & new_n1023_;
  assign new_n1042_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n459_ & new_n1023_;
  assign new_n1043_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n461_ & new_n1023_;
  assign new_n1044_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n463_ & new_n1023_;
  assign new_n1045_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n465_ & new_n1023_;
  assign new_n1046_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n467_ & new_n1023_;
  assign new_n1047_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n469_ & new_n1023_;
  assign new_n1048_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n471_ & new_n1023_;
  assign new_n1049_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n473_ & new_n1023_;
  assign new_n1050_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n475_ & new_n1023_;
  assign new_n1051_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n477_ & new_n1023_;
  assign new_n1052_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n479_ & new_n1023_;
  assign new_n1053_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n481_ & new_n1023_;
  assign new_n1054_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n483_ & new_n1023_;
  assign new_n1055_ = pi005 & new_n990_ & new_n924_ & new_n859_ & new_n957_ & new_n485_ & new_n1023_;
  assign new_n1056_ = ~pi005;
  assign new_n1057_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi111 & new_n1056_;
  assign new_n1058_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi112 & new_n1056_;
  assign new_n1059_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi113 & new_n1056_;
  assign new_n1060_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi114 & new_n1056_;
  assign new_n1061_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi115 & new_n1056_;
  assign new_n1062_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi116 & new_n1056_;
  assign new_n1063_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi117 & new_n1056_;
  assign new_n1064_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi118 & new_n1056_;
  assign new_n1065_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi119 & new_n1056_;
  assign new_n1066_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi120 & new_n1056_;
  assign new_n1067_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi121 & new_n1056_;
  assign new_n1068_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi122 & new_n1056_;
  assign new_n1069_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi123 & new_n1056_;
  assign new_n1070_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi124 & new_n1056_;
  assign new_n1071_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi125 & new_n1056_;
  assign new_n1072_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi110 & new_n1056_;
  assign new_n1073_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi107 & new_n1056_;
  assign new_n1074_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi108 & new_n1056_;
  assign new_n1075_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi109 & new_n1056_;
  assign new_n1076_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi106 & new_n1056_;
  assign new_n1077_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi104 & new_n1056_;
  assign new_n1078_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi105 & new_n1056_;
  assign new_n1079_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi103 & new_n1056_;
  assign new_n1080_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi097 & new_n1056_;
  assign new_n1081_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi098 & new_n1056_;
  assign new_n1082_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi099 & new_n1056_;
  assign new_n1083_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi100 & new_n1056_;
  assign new_n1084_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi101 & new_n1056_;
  assign new_n1085_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi102 & new_n1056_;
  assign new_n1086_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi094 & new_n1056_;
  assign new_n1087_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi096 & new_n1056_;
  assign new_n1088_ = new_n1355_ & pi095 & new_n1023_ & new_n957_ & new_n859_ & new_n924_ & new_n990_ & pi090 & new_n1056_;
  assign new_n1089_ = new_n1362_ & pi067;
  assign new_n1090_ = new_n1362_ & pi068;
  assign new_n1091_ = new_n1362_ & pi069;
  assign new_n1092_ = new_n1362_ & pi070;
  assign new_n1093_ = new_n1362_ & pi071;
  assign new_n1094_ = new_n1362_ & pi072;
  assign new_n1095_ = new_n1362_ & pi073;
  assign new_n1096_ = new_n1362_ & pi074;
  assign new_n1097_ = new_n1362_ & pi075;
  assign new_n1098_ = new_n1362_ & pi076;
  assign new_n1099_ = new_n1362_ & pi077;
  assign new_n1100_ = new_n1362_ & pi078;
  assign new_n1101_ = new_n1362_ & pi079;
  assign new_n1102_ = new_n1362_ & pi080;
  assign new_n1103_ = new_n1362_ & pi081;
  assign new_n1104_ = ~new_n1362_;
  assign new_n1105_ = new_n1104_ & pi067 & new_n1366_;
  assign po64 = new_n1136_ | new_n1089_ | new_n1105_ | new_n1152_ | new_n1154_;
  assign new_n1107_ = new_n1104_ & pi068 & new_n1366_;
  assign po65 = new_n1137_ | new_n1090_ | new_n1107_ | new_n1152_ | new_n1155_;
  assign new_n1109_ = new_n1104_ & pi069 & new_n1366_;
  assign po66 = new_n1138_ | new_n1091_ | new_n1109_ | new_n1152_ | new_n1156_;
  assign new_n1111_ = new_n1104_ & pi070 & new_n1366_;
  assign po67 = new_n1139_ | new_n1092_ | new_n1111_ | new_n1152_ | new_n1157_;
  assign new_n1113_ = new_n1104_ & pi071 & new_n1366_;
  assign po68 = new_n1140_ | new_n1093_ | new_n1113_ | new_n1152_ | new_n1158_;
  assign new_n1115_ = new_n1104_ & pi072 & new_n1366_;
  assign po69 = new_n1141_ | new_n1094_ | new_n1115_ | new_n1152_ | new_n1159_;
  assign new_n1117_ = new_n1104_ & pi073 & new_n1366_;
  assign po70 = new_n1142_ | new_n1095_ | new_n1117_ | new_n1152_ | new_n1160_;
  assign new_n1119_ = new_n1104_ & pi074 & new_n1366_;
  assign po71 = new_n1143_ | new_n1096_ | new_n1119_ | new_n1152_ | new_n1161_;
  assign new_n1121_ = new_n1104_ & pi075 & new_n1366_;
  assign po72 = new_n1144_ | new_n1097_ | new_n1121_ | new_n1152_ | new_n1162_;
  assign new_n1123_ = new_n1104_ & pi076 & new_n1366_;
  assign po73 = new_n1145_ | new_n1098_ | new_n1123_ | new_n1152_ | new_n1163_;
  assign new_n1125_ = new_n1104_ & pi077 & new_n1366_;
  assign po74 = new_n1146_ | new_n1099_ | new_n1125_ | new_n1152_ | new_n1164_;
  assign new_n1127_ = new_n1104_ & pi078 & new_n1366_;
  assign po75 = new_n1147_ | new_n1100_ | new_n1127_ | new_n1152_ | new_n1165_;
  assign new_n1129_ = new_n1104_ & pi079 & new_n1366_;
  assign po76 = new_n1148_ | new_n1101_ | new_n1129_ | new_n1152_ | new_n1166_;
  assign new_n1131_ = new_n1104_ & pi080 & new_n1366_;
  assign po77 = new_n1149_ | new_n1102_ | new_n1131_ | new_n1152_ | new_n1167_;
  assign new_n1133_ = new_n1104_ & pi081 & new_n1366_;
  assign po78 = new_n1150_ | new_n1103_ | new_n1133_ | new_n1152_ | new_n1168_;
  assign new_n1135_ = ~new_n1366_;
  assign new_n1136_ = pi005 & new_n1104_ & pi067 & new_n1135_;
  assign new_n1137_ = pi005 & new_n1104_ & pi068 & new_n1135_;
  assign new_n1138_ = pi005 & new_n1104_ & pi069 & new_n1135_;
  assign new_n1139_ = pi005 & new_n1104_ & pi070 & new_n1135_;
  assign new_n1140_ = pi005 & new_n1104_ & pi071 & new_n1135_;
  assign new_n1141_ = pi005 & new_n1104_ & pi072 & new_n1135_;
  assign new_n1142_ = pi005 & new_n1104_ & pi073 & new_n1135_;
  assign new_n1143_ = pi005 & new_n1104_ & pi074 & new_n1135_;
  assign new_n1144_ = pi005 & new_n1104_ & pi075 & new_n1135_;
  assign new_n1145_ = pi005 & new_n1104_ & pi076 & new_n1135_;
  assign new_n1146_ = pi005 & new_n1104_ & pi077 & new_n1135_;
  assign new_n1147_ = pi005 & new_n1104_ & pi078 & new_n1135_;
  assign new_n1148_ = pi005 & new_n1104_ & pi079 & new_n1135_;
  assign new_n1149_ = pi005 & new_n1104_ & pi080 & new_n1135_;
  assign new_n1150_ = pi005 & new_n1104_ & pi081 & new_n1135_;
  assign new_n1151_ = ~pi005;
  assign new_n1152_ = new_n1151_ & new_n1104_ & new_n1374_ & new_n1135_;
  assign new_n1153_ = ~new_n1374_;
  assign new_n1154_ = new_n1375_ & pi095 & new_n1151_ & new_n1104_ & new_n1135_ & pi108 & new_n1153_;
  assign new_n1155_ = new_n1375_ & pi095 & new_n1151_ & new_n1104_ & new_n1135_ & pi109 & new_n1153_;
  assign new_n1156_ = new_n1375_ & pi095 & new_n1151_ & new_n1104_ & new_n1135_ & pi106 & new_n1153_;
  assign new_n1157_ = new_n1375_ & pi095 & new_n1151_ & new_n1104_ & new_n1135_ & pi104 & new_n1153_;
  assign new_n1158_ = new_n1375_ & pi095 & new_n1151_ & new_n1104_ & new_n1135_ & pi105 & new_n1153_;
  assign new_n1159_ = new_n1375_ & pi095 & new_n1151_ & new_n1104_ & new_n1135_ & pi103 & new_n1153_;
  assign new_n1160_ = new_n1375_ & pi095 & new_n1151_ & new_n1104_ & new_n1135_ & pi097 & new_n1153_;
  assign new_n1161_ = new_n1375_ & pi095 & new_n1151_ & new_n1104_ & new_n1135_ & pi098 & new_n1153_;
  assign new_n1162_ = new_n1375_ & pi095 & new_n1151_ & new_n1104_ & new_n1135_ & pi099 & new_n1153_;
  assign new_n1163_ = new_n1375_ & pi095 & new_n1151_ & new_n1104_ & new_n1135_ & pi100 & new_n1153_;
  assign new_n1164_ = new_n1375_ & pi095 & new_n1151_ & new_n1104_ & new_n1135_ & pi101 & new_n1153_;
  assign new_n1165_ = new_n1375_ & pi095 & new_n1151_ & new_n1104_ & new_n1135_ & pi102 & new_n1153_;
  assign new_n1166_ = new_n1375_ & pi095 & new_n1151_ & new_n1104_ & new_n1135_ & pi094 & new_n1153_;
  assign new_n1167_ = new_n1375_ & pi095 & new_n1151_ & new_n1104_ & new_n1135_ & pi096 & new_n1153_;
  assign new_n1168_ = new_n1375_ & pi095 & new_n1151_ & new_n1104_ & new_n1135_ & pi090 & new_n1153_;
  assign new_n1169_ = new_n1379_ & pi126;
  assign new_n1170_ = ~new_n1379_;
  assign po79 = new_n1178_ | new_n1169_ | new_n1180_ | new_n1174_ | new_n1176_;
  assign new_n1172_ = ~new_n1381_;
  assign new_n1173_ = ~new_n1383_;
  assign new_n1174_ = pi005 & new_n1172_ & new_n1170_ & pi127 & new_n1173_;
  assign new_n1175_ = ~pi005;
  assign new_n1176_ = new_n1175_ & new_n1172_ & new_n1170_ & new_n1386_ & new_n1173_;
  assign new_n1177_ = ~new_n1386_;
  assign new_n1178_ = new_n1177_ & new_n1173_ & new_n1170_ & new_n1172_ & new_n1391_ & new_n1175_;
  assign new_n1179_ = ~new_n1391_;
  assign new_n1180_ = new_n1177_ & new_n1173_ & new_n1170_ & new_n1172_ & new_n1179_ & new_n1175_;
  assign new_n1181_ = new_n1394_ & pi128;
  assign new_n1182_ = ~new_n1394_;
  assign new_n1183_ = new_n1182_ & new_n1397_;
  assign po80 = new_n1186_ | new_n1181_ | new_n1183_;
  assign new_n1185_ = ~new_n1397_;
  assign new_n1186_ = pi005 & new_n1182_ & pi129 & new_n1185_;
  assign new_n1187_ = ~pi001;
  assign new_n1188_ = ~pi095;
  assign new_n1189_ = ~pi005;
  assign new_n1190_ = pi007 & new_n1188_ & new_n1189_ & new_n1187_;
  assign new_n1191_ = ~pi002;
  assign new_n1192_ = ~pi095;
  assign new_n1193_ = ~pi005;
  assign new_n1194_ = pi007 & new_n1191_ & new_n1193_ & new_n1192_;
  assign new_n1195_ = ~pi007;
  assign new_n1196_ = ~pi095;
  assign new_n1197_ = ~pi005;
  assign new_n1198_ = new_n1195_ & new_n1197_ & new_n1196_;
  assign new_n1199_ = ~pi005;
  assign new_n1200_ = new_n1199_ & pi095;
  assign new_n1201_ = ~pi130;
  assign new_n1202_ = ~pi008;
  assign new_n1203_ = ~pi095;
  assign new_n1204_ = new_n1201_ & new_n1202_ & pi002 & new_n1203_ & pi001;
  assign new_n1205_ = ~pi008;
  assign new_n1206_ = ~pi095;
  assign new_n1207_ = pi007 & new_n1206_ & new_n1205_;
  assign new_n1208_ = ~pi095;
  assign new_n1209_ = ~pi005;
  assign new_n1210_ = pi008 & new_n1209_ & new_n1208_;
  assign new_n1211_ = ~pi001;
  assign new_n1212_ = ~pi007;
  assign new_n1213_ = ~pi095;
  assign new_n1214_ = ~pi005;
  assign new_n1215_ = new_n1212_ & new_n1213_ & new_n1214_ & new_n1211_;
  assign new_n1216_ = ~pi002;
  assign new_n1217_ = ~pi007;
  assign new_n1218_ = ~pi095;
  assign new_n1219_ = ~pi005;
  assign new_n1220_ = new_n1217_ & new_n1216_ & new_n1219_ & new_n1218_;
  assign new_n1221_ = ~pi005;
  assign new_n1222_ = ~pi130;
  assign new_n1223_ = ~pi006;
  assign new_n1224_ = ~pi095;
  assign new_n1225_ = new_n1222_ & new_n1224_ & new_n1223_;
  assign new_n1226_ = ~pi095;
  assign new_n1227_ = new_n1226_ & pi007;
  assign new_n1228_ = ~pi005;
  assign new_n1229_ = ~pi130;
  assign new_n1230_ = ~pi095;
  assign new_n1231_ = new_n1230_ & new_n1229_;
  assign new_n1232_ = ~pi095;
  assign new_n1233_ = new_n1232_ & pi007;
  assign new_n1234_ = ~pi005;
  assign new_n1235_ = ~pi130;
  assign new_n1236_ = ~pi006;
  assign new_n1237_ = ~pi095;
  assign new_n1238_ = new_n1235_ & new_n1237_ & new_n1236_;
  assign new_n1239_ = ~pi095;
  assign new_n1240_ = new_n1239_ & pi007;
  assign new_n1241_ = ~pi005;
  assign new_n1242_ = ~pi001;
  assign new_n1243_ = ~pi130;
  assign new_n1244_ = ~pi095;
  assign new_n1245_ = new_n1243_ & new_n1244_ & new_n1242_;
  assign new_n1246_ = ~pi002;
  assign new_n1247_ = ~pi130;
  assign new_n1248_ = ~pi006;
  assign new_n1249_ = ~pi095;
  assign new_n1250_ = new_n1247_ & new_n1246_ & new_n1249_ & new_n1248_;
  assign new_n1251_ = ~pi130;
  assign new_n1252_ = ~pi095;
  assign new_n1253_ = pi000 & new_n1252_ & new_n1251_;
  assign new_n1254_ = ~pi095;
  assign new_n1255_ = new_n1254_ & pi007;
  assign new_n1256_ = ~pi005;
  assign new_n1257_ = new_n1256_ & pi095;
  assign new_n1258_ = ~pi000;
  assign new_n1259_ = ~pi130;
  assign new_n1260_ = ~pi007;
  assign new_n1261_ = ~pi095;
  assign new_n1262_ = ~pi005;
  assign new_n1263_ = ~pi001;
  assign new_n1264_ = ~pi130;
  assign new_n1265_ = ~pi006;
  assign new_n1266_ = ~pi095;
  assign new_n1267_ = new_n1264_ & new_n1265_ & new_n1266_ & new_n1263_;
  assign new_n1268_ = ~pi002;
  assign new_n1269_ = ~pi130;
  assign new_n1270_ = ~pi006;
  assign new_n1271_ = ~pi095;
  assign new_n1272_ = new_n1269_ & new_n1268_ & new_n1271_ & new_n1270_;
  assign new_n1273_ = ~pi130;
  assign new_n1274_ = ~pi095;
  assign new_n1275_ = pi000 & new_n1274_ & new_n1273_;
  assign new_n1276_ = ~pi095;
  assign new_n1277_ = new_n1276_ & pi007;
  assign new_n1278_ = ~pi005;
  assign new_n1279_ = new_n1278_ & pi095;
  assign new_n1280_ = ~pi000;
  assign new_n1281_ = ~pi130;
  assign new_n1282_ = ~pi007;
  assign new_n1283_ = ~pi095;
  assign new_n1284_ = ~pi005;
  assign new_n1285_ = ~pi001;
  assign new_n1286_ = ~pi002;
  assign new_n1287_ = ~pi130;
  assign new_n1288_ = ~pi095;
  assign new_n1289_ = new_n1287_ & new_n1286_ & new_n1288_ & new_n1285_;
  assign new_n1290_ = ~pi001;
  assign new_n1291_ = ~pi130;
  assign new_n1292_ = ~pi006;
  assign new_n1293_ = ~pi095;
  assign new_n1294_ = new_n1291_ & new_n1292_ & new_n1293_ & new_n1290_;
  assign new_n1295_ = ~pi002;
  assign new_n1296_ = ~pi130;
  assign new_n1297_ = ~pi006;
  assign new_n1298_ = ~pi095;
  assign new_n1299_ = new_n1296_ & new_n1295_ & new_n1298_ & new_n1297_;
  assign new_n1300_ = ~pi130;
  assign new_n1301_ = ~pi095;
  assign new_n1302_ = pi000 & new_n1301_ & new_n1300_;
  assign new_n1303_ = ~pi095;
  assign new_n1304_ = new_n1303_ & pi007;
  assign new_n1305_ = ~pi005;
  assign new_n1306_ = new_n1305_ & pi095;
  assign new_n1307_ = ~pi000;
  assign new_n1308_ = ~pi130;
  assign new_n1309_ = ~pi007;
  assign new_n1310_ = ~pi095;
  assign new_n1311_ = ~pi005;
  assign new_n1312_ = ~pi001;
  assign new_n1313_ = ~pi130;
  assign new_n1314_ = ~pi006;
  assign new_n1315_ = ~pi095;
  assign new_n1316_ = new_n1313_ & new_n1314_ & new_n1315_ & new_n1312_;
  assign new_n1317_ = ~pi002;
  assign new_n1318_ = ~pi130;
  assign new_n1319_ = ~pi006;
  assign new_n1320_ = ~pi095;
  assign new_n1321_ = new_n1318_ & new_n1317_ & new_n1320_ & new_n1319_;
  assign new_n1322_ = ~pi130;
  assign new_n1323_ = ~pi095;
  assign new_n1324_ = pi000 & new_n1323_ & new_n1322_;
  assign new_n1325_ = ~pi095;
  assign new_n1326_ = new_n1325_ & pi007;
  assign new_n1327_ = ~pi005;
  assign new_n1328_ = new_n1327_ & pi095;
  assign new_n1329_ = ~pi000;
  assign new_n1330_ = ~pi130;
  assign new_n1331_ = ~pi007;
  assign new_n1332_ = ~pi095;
  assign new_n1333_ = ~pi005;
  assign new_n1334_ = ~pi001;
  assign new_n1335_ = ~pi130;
  assign new_n1336_ = ~pi004;
  assign new_n1337_ = ~pi006;
  assign new_n1338_ = ~pi095;
  assign new_n1339_ = new_n1335_ & new_n1336_ & new_n1337_ & new_n1338_ & new_n1334_;
  assign new_n1340_ = ~pi001;
  assign new_n1341_ = ~pi095;
  assign new_n1342_ = ~pi131;
  assign new_n1343_ = pi004 & new_n1341_ & new_n1342_ & pi003 & new_n1340_;
  assign new_n1344_ = ~pi003;
  assign new_n1345_ = ~pi001;
  assign new_n1346_ = ~pi095;
  assign new_n1347_ = pi004 & new_n1346_ & new_n1344_ & new_n1345_;
  assign new_n1348_ = ~pi130;
  assign new_n1349_ = ~pi006;
  assign new_n1350_ = ~pi095;
  assign new_n1351_ = new_n1349_ & new_n1348_ & pi000 & pi002 & new_n1350_ & pi001;
  assign new_n1352_ = ~pi001;
  assign new_n1353_ = ~pi095;
  assign new_n1354_ = pi007 & new_n1353_ & new_n1352_;
  assign new_n1355_ = ~pi005;
  assign new_n1356_ = ~pi001;
  assign new_n1357_ = ~pi002;
  assign new_n1358_ = ~pi130;
  assign new_n1359_ = ~pi004;
  assign new_n1360_ = ~pi006;
  assign new_n1361_ = ~pi095;
  assign new_n1362_ = new_n1359_ & new_n1358_ & new_n1360_ & new_n1357_ & new_n1361_ & new_n1356_;
  assign new_n1363_ = ~pi001;
  assign new_n1364_ = ~pi002;
  assign new_n1365_ = ~pi095;
  assign new_n1366_ = pi007 & new_n1364_ & new_n1365_ & new_n1363_;
  assign new_n1367_ = ~pi001;
  assign new_n1368_ = ~pi002;
  assign new_n1369_ = ~pi007;
  assign new_n1370_ = ~pi095;
  assign new_n1371_ = ~pi005;
  assign new_n1372_ = ~pi131;
  assign new_n1373_ = ~pi132;
  assign new_n1374_ = new_n1369_ & new_n1370_ & pi004 & new_n1371_ & new_n1372_ & new_n1368_ & new_n1373_ & new_n1367_;
  assign new_n1375_ = ~pi005;
  assign new_n1376_ = ~pi008;
  assign new_n1377_ = ~pi095;
  assign new_n1378_ = ~pi005;
  assign new_n1379_ = pi007 & new_n1376_ & new_n1378_ & new_n1377_;
  assign new_n1380_ = ~pi005;
  assign new_n1381_ = new_n1380_ & pi095;
  assign new_n1382_ = ~pi005;
  assign new_n1383_ = pi002 & new_n1382_ & pi001;
  assign new_n1384_ = ~pi095;
  assign new_n1385_ = ~pi005;
  assign new_n1386_ = pi008 & new_n1385_ & new_n1384_;
  assign new_n1387_ = ~pi001;
  assign new_n1388_ = ~pi007;
  assign new_n1389_ = ~pi095;
  assign new_n1390_ = ~pi005;
  assign new_n1391_ = new_n1388_ & new_n1389_ & new_n1390_ & new_n1387_;
  assign new_n1392_ = ~pi095;
  assign new_n1393_ = ~pi005;
  assign new_n1394_ = pi007 & new_n1393_ & new_n1392_;
  assign new_n1395_ = ~pi095;
  assign new_n1396_ = ~pi005;
  assign new_n1397_ = new_n1395_ & pi002 & new_n1396_ & pi001;
endmodule


