// Benchmark "C7552.iscas" written by ABC on Thu Mar 19 13:02:36 2020

module C7552_iscas  ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107;
  wire new_n316_, new_n317_, new_n318_, new_n320_, new_n322_, new_n324_,
    new_n326_, new_n328_, new_n330_, new_n332_, new_n334_, new_n337_,
    new_n338_, new_n340_, new_n342_, new_n344_, new_n346_, new_n348_,
    new_n350_, new_n352_, new_n354_, new_n356_, new_n358_, new_n360_,
    new_n361_, new_n363_, new_n364_, new_n366_, new_n368_, new_n370_,
    new_n371_, new_n373_, new_n375_, new_n377_, new_n379_, new_n381_,
    new_n382_, new_n384_, new_n385_, new_n387_, new_n388_, new_n390_,
    new_n392_, new_n394_, new_n396_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n495_, new_n498_,
    new_n500_, new_n503_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_,
    new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_,
    new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_,
    new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_,
    new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_,
    new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_,
    new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_,
    new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_,
    new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_,
    new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_,
    new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_,
    new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_,
    new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_,
    new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_,
    new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_,
    new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_,
    new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_,
    new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_,
    new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_,
    new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_,
    new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_,
    new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_,
    new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_,
    new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_,
    new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_,
    new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_,
    new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_,
    new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_,
    new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_,
    new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_,
    new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_,
    new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_,
    new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_,
    new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_,
    new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_,
    new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_,
    new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_,
    new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_,
    new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_,
    new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_,
    new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_,
    new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_,
    new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_,
    new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_,
    new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_,
    new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_,
    new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_,
    new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_,
    new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_,
    new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_,
    new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_,
    new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_,
    new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_,
    new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_,
    new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_,
    new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_,
    new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_,
    new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_,
    new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_,
    new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_,
    new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_,
    new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_,
    new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_,
    new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_,
    new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_,
    new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_,
    new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_,
    new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_,
    new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_,
    new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_,
    new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_,
    new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_,
    new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_,
    new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_,
    new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_,
    new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_,
    new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_,
    new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_,
    new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_,
    new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_,
    new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_,
    new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_,
    new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_,
    new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_,
    new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_,
    new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_,
    new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_,
    new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_,
    new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_,
    new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_,
    new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_,
    new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_,
    new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_,
    new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_,
    new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_,
    new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_,
    new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_,
    new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_,
    new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_,
    new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_,
    new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_,
    new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_,
    new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_,
    new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_,
    new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_,
    new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_,
    new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_,
    new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_,
    new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_,
    new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_,
    new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_,
    new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_,
    new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_,
    new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_,
    new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_,
    new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_,
    new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_,
    new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_,
    new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_,
    new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_,
    new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_,
    new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_,
    new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_,
    new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_,
    new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_,
    new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_,
    new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_,
    new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_,
    new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_,
    new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_,
    new_n1847_, new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_,
    new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_,
    new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_,
    new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_,
    new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_,
    new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_,
    new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_,
    new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_,
    new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_,
    new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_,
    new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_,
    new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_,
    new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_,
    new_n1925_, new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_,
    new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_,
    new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_,
    new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_, new_n1948_,
    new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_,
    new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_,
    new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_,
    new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_,
    new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_,
    new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_,
    new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_,
    new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_,
    new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_,
    new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_,
    new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_,
    new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_,
    new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_,
    new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_,
    new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_,
    new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_,
    new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_,
    new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_,
    new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_,
    new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_,
    new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_,
    new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_,
    new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_,
    new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_,
    new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_,
    new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_,
    new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_,
    new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_,
    new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_,
    new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_,
    new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_,
    new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_,
    new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_,
    new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_,
    new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_,
    new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_,
    new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_, new_n2170_,
    new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_,
    new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_,
    new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_,
    new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_,
    new_n2195_, new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_,
    new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_,
    new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_,
    new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_,
    new_n2219_, new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_,
    new_n2225_, new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_,
    new_n2231_, new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_,
    new_n2237_, new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_,
    new_n2243_, new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_,
    new_n2249_, new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_,
    new_n2255_, new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_,
    new_n2261_, new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_,
    new_n2267_, new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_,
    new_n2273_, new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_,
    new_n2279_, new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_,
    new_n2285_, new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_,
    new_n2291_, new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_,
    new_n2297_, new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_,
    new_n2303_, new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_,
    new_n2309_, new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_,
    new_n2315_, new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_,
    new_n2321_, new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_,
    new_n2327_, new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_,
    new_n2333_, new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_,
    new_n2339_, new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_,
    new_n2345_, new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_,
    new_n2351_, new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_,
    new_n2357_, new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_,
    new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_,
    new_n2369_, new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_,
    new_n2375_, new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_,
    new_n2381_, new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_,
    new_n2387_, new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_,
    new_n2393_, new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_,
    new_n2399_, new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_,
    new_n2405_, new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_,
    new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_,
    new_n2417_, new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_,
    new_n2423_, new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_,
    new_n2429_, new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_,
    new_n2435_, new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_,
    new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_,
    new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_,
    new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_,
    new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_,
    new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_,
    new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_,
    new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_,
    new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_,
    new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_,
    new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_,
    new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_,
    new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_,
    new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_,
    new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_,
    new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_,
    new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_,
    new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_,
    new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_,
    new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_,
    new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_,
    new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_,
    new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_,
    new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_,
    new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_,
    new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_,
    new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_,
    new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_,
    new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_,
    new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_,
    new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_,
    new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_,
    new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_,
    new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_,
    new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_,
    new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_,
    new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_,
    new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_,
    new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_,
    new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_,
    new_n2675_, new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_,
    new_n2681_, new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_,
    new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_,
    new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_,
    new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_,
    new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_,
    new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_,
    new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_,
    new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_,
    new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_,
    new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_,
    new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_,
    new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_,
    new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_,
    new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_,
    new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_,
    new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_,
    new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_,
    new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_,
    new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_,
    new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_,
    new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_,
    new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_,
    new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_,
    new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_,
    new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_,
    new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_,
    new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_,
    new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_,
    new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_,
    new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_,
    new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_,
    new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_,
    new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_,
    new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_,
    new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_,
    new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_,
    new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_,
    new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_,
    new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_,
    new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_,
    new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_,
    new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_,
    new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_,
    new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_,
    new_n2945_, new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_,
    new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_,
    new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_,
    new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_,
    new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_,
    new_n2975_, new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_,
    new_n2981_, new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_,
    new_n2987_, new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_,
    new_n2993_, new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_,
    new_n2999_, new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_,
    new_n3005_, new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_,
    new_n3011_, new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_,
    new_n3017_, new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_,
    new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_,
    new_n3029_, new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_,
    new_n3035_, new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_,
    new_n3041_, new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_,
    new_n3047_, new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_,
    new_n3053_, new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_,
    new_n3059_, new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_,
    new_n3065_, new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_,
    new_n3071_, new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_,
    new_n3077_, new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_,
    new_n3083_, new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_,
    new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_,
    new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_,
    new_n3101_, new_n3102_, new_n3104_, new_n3105_, new_n3106_, new_n3107_,
    new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_,
    new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_,
    new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_,
    new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_,
    new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_,
    new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_,
    new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_,
    new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_,
    new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_,
    new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_,
    new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_,
    new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_,
    new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_,
    new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_,
    new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_,
    new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3205_, new_n3207_,
    new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_, new_n3213_,
    new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3220_, new_n3221_,
    new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_,
    new_n3228_, new_n3229_, new_n3232_, new_n3233_, new_n3234_, new_n3235_,
    new_n3236_, new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_,
    new_n3242_, new_n3243_, new_n3244_, new_n3245_, new_n3246_, new_n3247_,
    new_n3248_, new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_,
    new_n3254_, new_n3255_, new_n3256_, new_n3258_, new_n3259_, new_n3261_,
    new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_, new_n3267_,
    new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_, new_n3273_,
    new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_, new_n3279_,
    new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_, new_n3285_,
    new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_,
    new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_, new_n3297_,
    new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_, new_n3303_,
    new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_, new_n3309_,
    new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_, new_n3317_,
    new_n3318_, new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_,
    new_n3324_, new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_,
    new_n3330_, new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_,
    new_n3336_, new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_,
    new_n3342_, new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_,
    new_n3348_, new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_,
    new_n3354_, new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_,
    new_n3360_, new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_,
    new_n3366_, new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_,
    new_n3372_, new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_,
    new_n3378_, new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_,
    new_n3384_, new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_,
    new_n3390_, new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_,
    new_n3396_, new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_,
    new_n3402_, new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_,
    new_n3408_, new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_,
    new_n3414_, new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_,
    new_n3420_, new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_,
    new_n3426_, new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_,
    new_n3432_, new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_,
    new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_,
    new_n3444_, new_n3445_, new_n3446_, new_n3448_, new_n3449_, new_n3450_,
    new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3456_,
    new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3462_, new_n3463_,
    new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_,
    new_n3470_, new_n3471_, new_n3473_, new_n3474_, new_n3475_, new_n3476_,
    new_n3479_, new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_,
    new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_,
    new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3500_, new_n3501_,
    new_n3503_, new_n3504_, new_n3508_, new_n3509_, new_n3512_, new_n3513_,
    new_n3514_, new_n3515_, new_n3516_, new_n3518_, new_n3519_, new_n3522_,
    new_n3523_, new_n3524_, new_n3526_, new_n3528_, new_n3531_, new_n3532_,
    new_n3536_, new_n3537_, new_n3541_, new_n3542_, new_n3543_, new_n3544_,
    new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_,
    new_n3551_, new_n3552_, new_n3555_, new_n3556_, new_n3557_, new_n3562_,
    new_n3563_, new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_,
    new_n3569_, new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_,
    new_n3575_, new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_,
    new_n3581_, new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_,
    new_n3587_, new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_,
    new_n3593_, new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_,
    new_n3599_, new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_,
    new_n3605_, new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_,
    new_n3611_, new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_,
    new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_,
    new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_,
    new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_,
    new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_,
    new_n3641_, new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_,
    new_n3647_, new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_,
    new_n3653_, new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_,
    new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_,
    new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_,
    new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_,
    new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_,
    new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_,
    new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_,
    new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_,
    new_n3701_, new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_,
    new_n3707_, new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_,
    new_n3713_, new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_,
    new_n3719_, new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_,
    new_n3725_, new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_,
    new_n3731_, new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_,
    new_n3737_, new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_,
    new_n3743_, new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_,
    new_n3749_, new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_,
    new_n3755_, new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_,
    new_n3761_, new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_,
    new_n3767_, new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_,
    new_n3773_, new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_,
    new_n3779_, new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_,
    new_n3785_, new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_,
    new_n3791_, new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_,
    new_n3797_, new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_,
    new_n3803_, new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_,
    new_n3809_, new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_,
    new_n3815_, new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_,
    new_n3821_, new_n3822_, new_n3823_;
  assign new_n316_ = pi205;
  assign new_n317_ = pi205;
  assign new_n318_ = ~pi204;
  assign po036 = pi204;
  assign new_n320_ = ~pi203;
  assign po035 = pi203;
  assign new_n322_ = ~pi202;
  assign po034 = pi202;
  assign new_n324_ = ~pi201;
  assign po033 = pi201;
  assign new_n326_ = ~pi200;
  assign po032 = pi200;
  assign new_n328_ = ~pi199;
  assign po031 = pi199;
  assign new_n330_ = ~pi198;
  assign po030 = pi198;
  assign new_n332_ = ~pi197;
  assign po029 = pi197;
  assign new_n334_ = ~pi196;
  assign po040 = pi196;
  assign po028 = pi195;
  assign new_n337_ = ~pi195;
  assign new_n338_ = ~pi194;
  assign po027 = pi194;
  assign new_n340_ = ~pi193;
  assign po026 = pi193;
  assign new_n342_ = ~pi192;
  assign po025 = pi192;
  assign new_n344_ = ~pi191;
  assign po024 = pi191;
  assign new_n346_ = ~pi190;
  assign po023 = pi190;
  assign new_n348_ = ~pi189;
  assign po022 = pi189;
  assign new_n350_ = ~pi188;
  assign po021 = pi188;
  assign new_n352_ = ~pi187;
  assign po020 = pi187;
  assign new_n354_ = ~pi186;
  assign po019 = pi186;
  assign new_n356_ = ~pi185;
  assign po018 = pi185;
  assign new_n358_ = ~pi184;
  assign po017 = pi184;
  assign new_n360_ = ~pi184;
  assign new_n361_ = ~pi183;
  assign po016 = pi183;
  assign new_n363_ = ~pi183;
  assign new_n364_ = ~pi182;
  assign po015 = pi182;
  assign new_n366_ = ~pi181;
  assign po014 = pi181;
  assign new_n368_ = ~pi180;
  assign po013 = pi180;
  assign new_n370_ = ~pi180;
  assign new_n371_ = ~pi179;
  assign po012 = pi179;
  assign new_n373_ = ~pi178;
  assign po011 = pi178;
  assign new_n375_ = ~pi177;
  assign po010 = pi177;
  assign new_n377_ = ~pi176;
  assign po039 = pi176;
  assign new_n379_ = ~pi175;
  assign po009 = pi175;
  assign new_n381_ = ~pi174;
  assign new_n382_ = ~pi173;
  assign po008 = pi173;
  assign new_n384_ = ~pi206 | ~pi173;
  assign new_n385_ = ~pi172;
  assign po007 = pi172;
  assign new_n387_ = pi206 & pi172;
  assign new_n388_ = ~pi171;
  assign po006 = pi171;
  assign new_n390_ = ~pi170;
  assign po005 = pi170;
  assign new_n392_ = ~pi169;
  assign po004 = pi169;
  assign new_n394_ = ~pi168;
  assign po038 = pi168;
  assign new_n396_ = ~pi167;
  assign po003 = pi167;
  assign new_n398_ = ~pi166;
  assign new_n399_ = pi109 & pi108 & pi106 & pi105;
  assign new_n400_ = pi122 & pi111 & pi085 & pi095;
  assign new_n401_ = pi153 & pi141 & pi133 & pi075;
  assign new_n402_ = pi163 & pi151 & pi073 & pi107;
  assign new_n403_ = pi067 & pi066;
  assign new_n404_ = pi053;
  assign new_n405_ = ~pi053;
  assign new_n406_ = ~pi020;
  assign new_n407_ = pi011;
  assign new_n408_ = pi011;
  assign new_n409_ = pi005;
  assign new_n410_ = pi005;
  assign new_n411_ = ~pi005;
  assign new_n412_ = pi005;
  assign po037 = ~pi004;
  assign new_n414_ = pi004;
  assign new_n415_ = ~pi003 | ~pi002;
  assign new_n416_ = ~pi003 | ~pi002;
  assign new_n417_ = ~pi001;
  assign new_n418_ = ~pi001;
  assign new_n419_ = ~pi001;
  assign new_n420_ = pi000;
  assign po002 = pi000;
  assign po001 = pi000;
  assign new_n423_ = ~pi206 | ~new_n381_;
  assign new_n424_ = pi206 & new_n398_;
  assign new_n425_ = ~new_n316_;
  assign new_n426_ = ~new_n317_;
  assign new_n427_ = new_n318_;
  assign new_n428_ = new_n318_;
  assign new_n429_ = new_n320_;
  assign new_n430_ = new_n320_;
  assign new_n431_ = new_n322_;
  assign new_n432_ = new_n322_;
  assign new_n433_ = new_n324_;
  assign new_n434_ = new_n324_;
  assign new_n435_ = new_n326_;
  assign new_n436_ = new_n326_;
  assign new_n437_ = new_n328_;
  assign new_n438_ = new_n328_;
  assign new_n439_ = new_n330_;
  assign new_n440_ = new_n330_;
  assign new_n441_ = new_n332_;
  assign new_n442_ = new_n332_;
  assign new_n443_ = new_n334_;
  assign new_n444_ = new_n334_;
  assign new_n445_ = new_n338_;
  assign new_n446_ = new_n338_;
  assign new_n447_ = new_n340_;
  assign new_n448_ = new_n340_;
  assign new_n449_ = new_n342_;
  assign new_n450_ = new_n342_;
  assign new_n451_ = new_n344_;
  assign new_n452_ = new_n344_;
  assign new_n453_ = new_n346_;
  assign new_n454_ = new_n346_;
  assign new_n455_ = new_n348_;
  assign new_n456_ = new_n348_;
  assign new_n457_ = new_n350_;
  assign new_n458_ = new_n350_;
  assign new_n459_ = new_n352_;
  assign new_n460_ = new_n352_;
  assign new_n461_ = new_n360_;
  assign new_n462_ = new_n360_;
  assign new_n463_ = new_n363_;
  assign new_n464_ = new_n363_;
  assign new_n465_ = new_n364_;
  assign new_n466_ = new_n364_;
  assign new_n467_ = new_n366_;
  assign new_n468_ = new_n366_;
  assign new_n469_ = new_n370_;
  assign new_n470_ = new_n370_;
  assign new_n471_ = new_n371_;
  assign new_n472_ = new_n371_;
  assign new_n473_ = new_n373_;
  assign new_n474_ = new_n373_;
  assign new_n475_ = new_n375_;
  assign new_n476_ = new_n375_;
  assign new_n477_ = new_n377_;
  assign new_n478_ = new_n377_;
  assign new_n479_ = new_n384_ & new_n408_;
  assign new_n480_ = new_n384_ & new_n408_;
  assign new_n481_ = new_n384_;
  assign new_n482_ = new_n384_;
  assign new_n483_ = ~new_n387_;
  assign new_n484_ = new_n388_;
  assign new_n485_ = new_n388_;
  assign new_n486_ = new_n390_;
  assign new_n487_ = new_n390_;
  assign new_n488_ = new_n392_;
  assign new_n489_ = new_n392_;
  assign new_n490_ = new_n394_;
  assign new_n491_ = new_n394_;
  assign po050 = ~pi165 | ~new_n417_;
  assign po048 = ~pi165 | ~new_n417_;
  assign po044 = ~new_n399_;
  assign new_n495_ = new_n399_ & new_n400_;
  assign po045 = ~new_n400_;
  assign po043 = ~new_n401_;
  assign new_n498_ = new_n402_ & new_n401_;
  assign po042 = ~new_n402_;
  assign new_n500_ = new_n403_ & new_n418_;
  assign po051 = ~new_n403_ | ~new_n418_;
  assign po047 = new_n404_;
  assign new_n503_ = ~new_n404_;
  assign po041 = ~new_n406_ | ~new_n419_;
  assign new_n505_ = new_n407_;
  assign new_n506_ = new_n407_;
  assign new_n507_ = new_n408_;
  assign new_n508_ = new_n408_;
  assign new_n509_ = new_n408_;
  assign new_n510_ = new_n408_;
  assign new_n511_ = new_n409_;
  assign new_n512_ = new_n409_;
  assign new_n513_ = new_n409_;
  assign new_n514_ = new_n409_;
  assign new_n515_ = ~new_n409_;
  assign new_n516_ = new_n410_;
  assign new_n517_ = new_n410_;
  assign new_n518_ = new_n410_;
  assign new_n519_ = new_n410_;
  assign new_n520_ = ~new_n410_;
  assign new_n521_ = new_n411_;
  assign new_n522_ = new_n411_;
  assign new_n523_ = new_n412_;
  assign new_n524_ = new_n412_;
  assign new_n525_ = new_n412_;
  assign new_n526_ = new_n412_;
  assign new_n527_ = ~new_n412_;
  assign po049 = ~new_n414_;
  assign po052 = ~new_n414_;
  assign new_n530_ = new_n415_;
  assign new_n531_ = new_n415_;
  assign new_n532_ = new_n415_;
  assign new_n533_ = new_n416_;
  assign new_n534_ = new_n416_;
  assign new_n535_ = new_n416_;
  assign new_n536_ = new_n420_;
  assign po046 = new_n420_;
  assign new_n538_ = new_n423_;
  assign new_n539_ = ~new_n424_;
  assign new_n540_ = ~new_n427_;
  assign new_n541_ = ~new_n428_;
  assign new_n542_ = ~new_n429_;
  assign new_n543_ = ~new_n430_;
  assign new_n544_ = ~new_n431_;
  assign new_n545_ = ~new_n432_;
  assign new_n546_ = ~new_n433_;
  assign new_n547_ = ~new_n434_;
  assign new_n548_ = ~new_n435_;
  assign new_n549_ = ~new_n436_;
  assign new_n550_ = ~new_n437_;
  assign new_n551_ = ~new_n438_;
  assign new_n552_ = ~new_n439_;
  assign new_n553_ = ~new_n440_;
  assign new_n554_ = ~new_n441_;
  assign new_n555_ = ~new_n442_;
  assign new_n556_ = ~new_n443_;
  assign new_n557_ = ~new_n444_;
  assign new_n558_ = ~new_n445_;
  assign new_n559_ = ~new_n446_;
  assign new_n560_ = ~new_n447_;
  assign new_n561_ = ~new_n448_;
  assign new_n562_ = ~new_n449_;
  assign new_n563_ = ~new_n450_;
  assign new_n564_ = ~new_n451_;
  assign new_n565_ = ~new_n452_;
  assign new_n566_ = ~new_n453_;
  assign new_n567_ = ~new_n454_;
  assign new_n568_ = ~new_n455_;
  assign new_n569_ = ~new_n456_;
  assign new_n570_ = ~new_n457_;
  assign new_n571_ = ~new_n458_;
  assign new_n572_ = ~new_n459_;
  assign new_n573_ = ~new_n460_;
  assign new_n574_ = new_n358_ & new_n519_;
  assign new_n575_ = ~new_n461_;
  assign new_n576_ = ~new_n462_;
  assign new_n577_ = new_n361_ & new_n519_;
  assign new_n578_ = ~new_n463_;
  assign new_n579_ = ~new_n464_;
  assign new_n580_ = new_n364_ & new_n519_;
  assign new_n581_ = ~new_n465_;
  assign new_n582_ = ~new_n466_;
  assign new_n583_ = ~new_n467_;
  assign new_n584_ = ~new_n468_;
  assign new_n585_ = new_n366_ & new_n519_;
  assign new_n586_ = new_n368_ & new_n519_;
  assign new_n587_ = ~new_n469_;
  assign new_n588_ = ~new_n470_;
  assign new_n589_ = ~new_n471_;
  assign new_n590_ = ~new_n472_;
  assign new_n591_ = new_n371_ & new_n518_;
  assign new_n592_ = new_n373_ & new_n518_;
  assign new_n593_ = ~new_n473_;
  assign new_n594_ = ~new_n474_;
  assign new_n595_ = ~new_n475_;
  assign new_n596_ = ~new_n476_;
  assign new_n597_ = new_n375_ & new_n518_;
  assign new_n598_ = ~new_n477_;
  assign new_n599_ = new_n377_ & new_n518_;
  assign new_n600_ = ~new_n478_;
  assign new_n601_ = new_n379_ & new_n518_;
  assign new_n602_ = new_n382_ & new_n517_;
  assign new_n603_ = ~new_n481_;
  assign new_n604_ = ~new_n482_;
  assign new_n605_ = new_n385_ & new_n517_;
  assign new_n606_ = new_n483_;
  assign new_n607_ = new_n483_;
  assign new_n608_ = new_n388_ & new_n517_;
  assign new_n609_ = ~new_n484_;
  assign new_n610_ = ~new_n485_;
  assign new_n611_ = ~new_n486_;
  assign new_n612_ = ~new_n487_;
  assign new_n613_ = new_n390_ & new_n516_;
  assign new_n614_ = ~new_n488_;
  assign new_n615_ = new_n392_ & new_n516_;
  assign new_n616_ = ~new_n489_;
  assign new_n617_ = ~new_n490_;
  assign new_n618_ = new_n394_ & new_n516_;
  assign new_n619_ = ~new_n491_;
  assign new_n620_ = new_n396_ & new_n516_;
  assign new_n621_ = pi139 & new_n525_;
  assign new_n622_ = pi138 & new_n525_;
  assign new_n623_ = pi137 & new_n525_;
  assign new_n624_ = pi136 & new_n526_;
  assign new_n625_ = pi135 & new_n526_;
  assign new_n626_ = pi134 & new_n526_;
  assign new_n627_ = pi132 & new_n525_;
  assign new_n628_ = pi104 & new_n514_;
  assign new_n629_ = pi103 & new_n514_;
  assign new_n630_ = pi102 & new_n514_;
  assign new_n631_ = pi101 & new_n514_;
  assign new_n632_ = pi100 & new_n513_;
  assign new_n633_ = pi099 & new_n513_;
  assign new_n634_ = pi098 & new_n513_;
  assign new_n635_ = pi097 & new_n513_;
  assign new_n636_ = pi096 & new_n513_;
  assign new_n637_ = pi094 & new_n514_;
  assign new_n638_ = pi093 & new_n511_;
  assign new_n639_ = pi092 & new_n511_;
  assign new_n640_ = pi091 & new_n511_;
  assign new_n641_ = pi090 & new_n511_;
  assign new_n642_ = pi089 & new_n512_;
  assign new_n643_ = pi088 & new_n512_;
  assign new_n644_ = pi087 & new_n512_;
  assign po055 = pi086 & new_n536_;
  assign new_n646_ = pi084 & new_n524_;
  assign new_n647_ = pi083 & new_n524_;
  assign new_n648_ = pi082 & new_n524_;
  assign new_n649_ = pi081 & new_n524_;
  assign new_n650_ = pi080 & new_n523_;
  assign new_n651_ = pi079 & new_n523_;
  assign new_n652_ = pi078 & new_n523_;
  assign new_n653_ = pi077 & new_n523_;
  assign new_n654_ = pi076 & new_n523_;
  assign new_n655_ = pi074 & new_n524_;
  assign po053 = ~new_n500_;
  assign new_n657_ = new_n503_;
  assign new_n658_ = new_n503_;
  assign new_n659_ = new_n405_ & new_n516_;
  assign new_n660_ = pi029 & new_n521_;
  assign new_n661_ = pi015 & new_n521_;
  assign new_n662_ = pi014 & new_n521_;
  assign new_n663_ = pi013 & new_n522_;
  assign new_n664_ = pi012 & new_n522_;
  assign new_n665_ = ~new_n505_;
  assign new_n666_ = new_n423_ & new_n407_;
  assign new_n667_ = ~new_n506_;
  assign new_n668_ = new_n483_ & new_n408_;
  assign new_n669_ = new_n408_ & new_n483_;
  assign new_n670_ = ~new_n408_ & ~new_n483_;
  assign new_n671_ = ~new_n507_;
  assign new_n672_ = ~new_n508_;
  assign new_n673_ = ~new_n483_ & ~new_n408_;
  assign new_n674_ = ~new_n509_;
  assign new_n675_ = ~new_n510_;
  assign new_n676_ = pi010 & new_n521_;
  assign new_n677_ = pi009 & new_n521_;
  assign new_n678_ = pi008 & new_n522_;
  assign new_n679_ = pi007 & new_n522_;
  assign new_n680_ = pi006 & new_n522_;
  assign new_n681_ = ~new_n511_;
  assign new_n682_ = ~new_n512_;
  assign new_n683_ = ~new_n513_;
  assign new_n684_ = ~new_n514_;
  assign new_n685_ = new_n515_;
  assign new_n686_ = new_n515_;
  assign new_n687_ = ~new_n516_;
  assign new_n688_ = ~new_n517_;
  assign new_n689_ = ~new_n518_;
  assign new_n690_ = ~new_n519_;
  assign new_n691_ = new_n520_;
  assign new_n692_ = new_n520_;
  assign new_n693_ = new_n520_;
  assign new_n694_ = new_n520_;
  assign new_n695_ = ~new_n521_;
  assign new_n696_ = ~new_n522_;
  assign new_n697_ = ~new_n523_;
  assign new_n698_ = ~new_n524_;
  assign new_n699_ = ~new_n525_;
  assign new_n700_ = ~new_n526_;
  assign new_n701_ = new_n527_;
  assign new_n702_ = new_n527_;
  assign new_n703_ = new_n527_;
  assign new_n704_ = new_n527_;
  assign po054 = new_n536_;
  assign new_n706_ = ~new_n538_ | ~new_n667_;
  assign new_n707_ = ~new_n538_;
  assign new_n708_ = new_n539_;
  assign new_n709_ = new_n354_ & new_n688_;
  assign new_n710_ = pi174 & new_n688_;
  assign new_n711_ = ~new_n481_ | ~new_n672_;
  assign new_n712_ = ~new_n482_ | ~new_n675_;
  assign new_n713_ = ~new_n606_ | ~new_n674_;
  assign new_n714_ = ~new_n606_;
  assign new_n715_ = ~new_n607_ | ~new_n671_;
  assign new_n716_ = ~new_n607_;
  assign new_n717_ = pi166 & new_n688_;
  assign new_n718_ = new_n699_ | new_n621_;
  assign new_n719_ = new_n699_ | new_n622_;
  assign new_n720_ = new_n699_ | new_n623_;
  assign new_n721_ = new_n700_ | new_n624_;
  assign new_n722_ = new_n700_ | new_n625_;
  assign new_n723_ = new_n700_ | new_n626_;
  assign new_n724_ = new_n699_ | new_n627_;
  assign new_n725_ = pi131 & new_n696_;
  assign new_n726_ = pi130 & new_n696_;
  assign new_n727_ = pi129 & new_n696_;
  assign new_n728_ = pi128 & new_n696_;
  assign new_n729_ = pi121 & new_n696_;
  assign new_n730_ = pi116 & new_n695_;
  assign new_n731_ = pi115 & new_n695_;
  assign new_n732_ = pi114 & new_n695_;
  assign new_n733_ = pi113 & new_n695_;
  assign new_n734_ = pi112 & new_n695_;
  assign new_n735_ = new_n683_ | new_n632_;
  assign new_n736_ = new_n683_ | new_n633_;
  assign new_n737_ = new_n683_ | new_n634_;
  assign new_n738_ = new_n683_ | new_n635_;
  assign new_n739_ = new_n683_ | new_n636_;
  assign new_n740_ = new_n681_ | new_n638_;
  assign new_n741_ = new_n681_ | new_n639_;
  assign new_n742_ = new_n681_ | new_n640_;
  assign new_n743_ = new_n681_ | new_n641_;
  assign new_n744_ = new_n682_ | new_n642_;
  assign new_n745_ = new_n682_ | new_n643_;
  assign new_n746_ = new_n682_ | new_n644_;
  assign new_n747_ = new_n697_ | new_n650_;
  assign new_n748_ = new_n697_ | new_n651_;
  assign new_n749_ = new_n697_ | new_n652_;
  assign new_n750_ = new_n697_ | new_n653_;
  assign new_n751_ = new_n697_ | new_n654_;
  assign new_n752_ = pi072 & new_n698_;
  assign new_n753_ = pi072 & new_n684_;
  assign new_n754_ = pi071 & new_n698_;
  assign new_n755_ = pi071 & new_n684_;
  assign new_n756_ = pi070 & new_n684_;
  assign new_n757_ = pi070 & new_n698_;
  assign new_n758_ = pi069 & new_n698_;
  assign new_n759_ = pi069 & new_n684_;
  assign new_n760_ = pi068 & new_n698_;
  assign new_n761_ = pi068 & new_n684_;
  assign new_n762_ = pi065 & new_n685_;
  assign new_n763_ = pi065 & new_n701_;
  assign new_n764_ = pi064 & new_n701_;
  assign new_n765_ = pi064 & new_n685_;
  assign new_n766_ = pi063 & new_n701_;
  assign new_n767_ = pi063 & new_n685_;
  assign new_n768_ = pi062 & new_n702_;
  assign new_n769_ = pi062 & new_n686_;
  assign new_n770_ = pi061 & new_n686_;
  assign new_n771_ = pi061 & new_n702_;
  assign new_n772_ = pi060 & new_n686_;
  assign new_n773_ = pi060 & new_n702_;
  assign new_n774_ = pi059 & new_n687_;
  assign new_n775_ = pi058 & new_n687_;
  assign new_n776_ = pi057 & new_n687_;
  assign new_n777_ = pi056 & new_n687_;
  assign new_n778_ = pi055 & new_n690_;
  assign new_n779_ = pi054 & new_n690_;
  assign new_n780_ = ~new_n657_;
  assign new_n781_ = ~new_n658_;
  assign new_n782_ = pi052 & new_n685_;
  assign new_n783_ = pi052 & new_n701_;
  assign new_n784_ = pi051 & new_n701_;
  assign new_n785_ = pi051 & new_n685_;
  assign new_n786_ = pi050 & new_n702_;
  assign new_n787_ = pi050 & new_n686_;
  assign new_n788_ = pi049 & new_n702_;
  assign new_n789_ = pi049 & new_n686_;
  assign new_n790_ = pi047 & new_n688_;
  assign new_n791_ = pi046 & new_n687_;
  assign new_n792_ = pi045 & new_n690_;
  assign new_n793_ = pi044 & new_n689_;
  assign new_n794_ = pi043 & new_n689_;
  assign new_n795_ = pi042 & new_n689_;
  assign new_n796_ = pi041 & new_n689_;
  assign new_n797_ = pi040 & new_n693_;
  assign new_n798_ = pi039 & new_n694_;
  assign new_n799_ = pi038 & new_n694_;
  assign new_n800_ = pi037 & new_n693_;
  assign new_n801_ = pi036 & new_n693_;
  assign new_n802_ = pi035 & new_n691_;
  assign new_n803_ = pi034 & new_n691_;
  assign new_n804_ = pi033 & new_n691_;
  assign new_n805_ = pi032 & new_n692_;
  assign new_n806_ = pi031 & new_n691_;
  assign new_n807_ = pi031 & new_n688_;
  assign new_n808_ = pi030 & new_n691_;
  assign new_n809_ = pi029 & new_n704_;
  assign new_n810_ = pi028 & new_n689_;
  assign new_n811_ = pi027 & new_n690_;
  assign new_n812_ = pi026 & new_n690_;
  assign new_n813_ = pi025 & new_n694_;
  assign new_n814_ = pi024 & new_n694_;
  assign new_n815_ = pi023 & new_n694_;
  assign new_n816_ = pi022 & new_n693_;
  assign new_n817_ = pi021 & new_n693_;
  assign new_n818_ = pi019 & new_n692_;
  assign new_n819_ = pi018 & new_n692_;
  assign new_n820_ = pi017 & new_n692_;
  assign new_n821_ = pi016 & new_n692_;
  assign new_n822_ = pi015 & new_n704_;
  assign new_n823_ = pi014 & new_n704_;
  assign new_n824_ = pi013 & new_n703_;
  assign new_n825_ = pi012 & new_n703_;
  assign new_n826_ = new_n539_ & new_n407_;
  assign new_n827_ = new_n668_;
  assign new_n828_ = new_n669_;
  assign new_n829_ = ~new_n670_;
  assign new_n830_ = ~new_n508_ | ~new_n603_;
  assign new_n831_ = ~new_n673_;
  assign new_n832_ = ~new_n510_ | ~new_n604_;
  assign new_n833_ = pi010 & new_n704_;
  assign new_n834_ = pi009 & new_n704_;
  assign new_n835_ = pi008 & new_n703_;
  assign new_n836_ = pi007 & new_n703_;
  assign new_n837_ = pi006 & new_n703_;
  assign new_n838_ = new_n681_ | new_n511_;
  assign new_n839_ = ~new_n685_;
  assign new_n840_ = ~new_n686_;
  assign new_n841_ = ~new_n691_;
  assign new_n842_ = ~new_n692_;
  assign new_n843_ = ~new_n693_;
  assign new_n844_ = ~new_n694_;
  assign new_n845_ = new_n699_ | new_n525_;
  assign new_n846_ = ~new_n701_;
  assign new_n847_ = ~new_n702_;
  assign new_n848_ = ~new_n703_;
  assign new_n849_ = ~new_n704_;
  assign new_n850_ = ~new_n708_;
  assign new_n851_ = new_n318_ & new_n844_;
  assign new_n852_ = new_n320_ & new_n844_;
  assign new_n853_ = new_n322_ & new_n844_;
  assign new_n854_ = new_n324_ & new_n844_;
  assign new_n855_ = new_n326_ & new_n844_;
  assign new_n856_ = new_n328_ & new_n843_;
  assign new_n857_ = new_n330_ & new_n843_;
  assign new_n858_ = new_n332_ & new_n843_;
  assign new_n859_ = new_n334_ & new_n843_;
  assign new_n860_ = new_n337_ & new_n843_;
  assign new_n861_ = new_n338_ & new_n842_;
  assign new_n862_ = new_n340_ & new_n842_;
  assign new_n863_ = new_n342_ & new_n842_;
  assign new_n864_ = new_n344_ & new_n842_;
  assign new_n865_ = new_n346_ & new_n842_;
  assign new_n866_ = new_n348_ & new_n841_;
  assign new_n867_ = new_n350_ & new_n841_;
  assign new_n868_ = new_n352_ & new_n841_;
  assign new_n869_ = new_n354_ & new_n841_;
  assign new_n870_ = new_n356_ & new_n841_;
  assign new_n871_ = new_n778_ | new_n574_;
  assign new_n872_ = new_n779_ | new_n577_;
  assign new_n873_ = new_n792_ | new_n580_;
  assign new_n874_ = new_n812_ | new_n585_;
  assign new_n875_ = new_n811_ | new_n586_;
  assign new_n876_ = new_n793_ | new_n591_;
  assign new_n877_ = new_n794_ | new_n592_;
  assign new_n878_ = new_n795_ | new_n597_;
  assign new_n879_ = new_n810_ | new_n599_;
  assign new_n880_ = new_n796_ | new_n601_;
  assign new_n881_ = new_n710_ | new_n602_;
  assign new_n882_ = ~new_n830_ | ~new_n711_;
  assign new_n883_ = ~new_n832_ | ~new_n712_;
  assign new_n884_ = new_n717_ | new_n605_;
  assign new_n885_ = new_n790_ | new_n608_;
  assign new_n886_ = new_n776_ | new_n613_;
  assign new_n887_ = new_n777_ | new_n615_;
  assign new_n888_ = new_n775_ | new_n618_;
  assign new_n889_ = new_n774_ | new_n620_;
  assign new_n890_ = pi162 & new_n848_;
  assign new_n891_ = pi161 & new_n848_;
  assign new_n892_ = pi160 & new_n848_;
  assign new_n893_ = pi159 & new_n848_;
  assign new_n894_ = pi158 & new_n846_;
  assign new_n895_ = pi157 & new_n846_;
  assign new_n896_ = pi156 & new_n846_;
  assign new_n897_ = pi155 & new_n846_;
  assign new_n898_ = pi154 & new_n846_;
  assign new_n899_ = pi152 & new_n848_;
  assign new_n900_ = pi150 & new_n847_;
  assign new_n901_ = pi149 & new_n847_;
  assign new_n902_ = pi148 & new_n847_;
  assign new_n903_ = pi147 & new_n847_;
  assign new_n904_ = pi146 & new_n849_;
  assign new_n905_ = pi145 & new_n849_;
  assign new_n906_ = pi144 & new_n849_;
  assign new_n907_ = pi143 & new_n849_;
  assign new_n908_ = pi142 & new_n849_;
  assign new_n909_ = pi140 & new_n847_;
  assign new_n910_ = pi127 & new_n839_;
  assign new_n911_ = pi126 & new_n839_;
  assign new_n912_ = pi125 & new_n839_;
  assign new_n913_ = pi124 & new_n839_;
  assign new_n914_ = pi123 & new_n839_;
  assign new_n915_ = pi120 & new_n840_;
  assign new_n916_ = pi119 & new_n840_;
  assign new_n917_ = pi118 & new_n840_;
  assign new_n918_ = pi117 & new_n840_;
  assign new_n919_ = pi110 & new_n840_;
  assign new_n920_ = new_n756_ | new_n628_;
  assign new_n921_ = new_n759_ | new_n629_;
  assign new_n922_ = new_n755_ | new_n630_;
  assign new_n923_ = new_n761_ | new_n631_;
  assign new_n924_ = new_n753_ | new_n637_;
  assign new_n925_ = new_n757_ | new_n646_;
  assign new_n926_ = new_n758_ | new_n647_;
  assign new_n927_ = new_n754_ | new_n648_;
  assign new_n928_ = new_n760_ | new_n649_;
  assign new_n929_ = new_n752_ | new_n655_;
  assign new_n930_ = new_n791_ | new_n659_;
  assign new_n931_ = new_n734_ | new_n660_;
  assign new_n932_ = new_n733_ | new_n661_;
  assign new_n933_ = new_n730_ | new_n662_;
  assign new_n934_ = new_n725_ | new_n663_;
  assign new_n935_ = new_n729_ | new_n664_;
  assign new_n936_ = ~new_n708_ | ~new_n665_;
  assign new_n937_ = ~new_n506_ | ~new_n707_;
  assign new_n938_ = ~new_n827_;
  assign new_n939_ = ~new_n828_;
  assign new_n940_ = ~new_n507_ | ~new_n716_;
  assign new_n941_ = ~new_n509_ | ~new_n714_;
  assign new_n942_ = new_n731_ | new_n676_;
  assign new_n943_ = new_n732_ | new_n677_;
  assign new_n944_ = new_n726_ | new_n678_;
  assign new_n945_ = new_n727_ | new_n679_;
  assign new_n946_ = new_n728_ | new_n680_;
  assign new_n947_ = new_n807_ | new_n517_;
  assign new_n948_ = new_n709_ | new_n517_;
  assign new_n949_ = new_n740_ & new_n530_;
  assign new_n950_ = new_n743_ & new_n530_;
  assign new_n951_ = new_n742_ & new_n530_;
  assign new_n952_ = new_n741_ & new_n530_;
  assign new_n953_ = new_n838_ & new_n530_;
  assign new_n954_ = new_n746_ & new_n531_;
  assign new_n955_ = new_n745_ & new_n531_;
  assign new_n956_ = new_n744_ & new_n531_;
  assign new_n957_ = new_n739_ & new_n532_;
  assign new_n958_ = new_n738_ & new_n532_;
  assign new_n959_ = new_n737_ & new_n532_;
  assign new_n960_ = new_n736_ & new_n532_;
  assign new_n961_ = new_n735_ & new_n532_;
  assign new_n962_ = new_n749_ & new_n533_;
  assign new_n963_ = new_n748_ & new_n533_;
  assign new_n964_ = new_n747_ & new_n533_;
  assign new_n965_ = new_n751_ & new_n533_;
  assign new_n966_ = new_n750_ & new_n533_;
  assign new_n967_ = new_n720_ & new_n534_;
  assign new_n968_ = new_n719_ & new_n534_;
  assign new_n969_ = new_n718_ & new_n534_;
  assign new_n970_ = new_n724_ & new_n534_;
  assign new_n971_ = new_n845_ & new_n534_;
  assign new_n972_ = new_n723_ & new_n535_;
  assign new_n973_ = new_n722_ & new_n535_;
  assign new_n974_ = new_n721_ & new_n535_;
  assign new_n975_ = ~new_n937_ | ~new_n706_;
  assign new_n976_ = new_n871_ & new_n957_;
  assign new_n977_ = new_n871_;
  assign new_n978_ = new_n871_;
  assign new_n979_ = new_n360_ & new_n965_;
  assign new_n980_ = new_n360_ & new_n965_;
  assign new_n981_ = new_n872_ & new_n958_;
  assign new_n982_ = new_n872_;
  assign new_n983_ = new_n872_;
  assign new_n984_ = new_n363_ & new_n966_;
  assign new_n985_ = new_n363_ & new_n966_;
  assign new_n986_ = new_n364_ & new_n962_;
  assign new_n987_ = new_n364_ & new_n962_;
  assign new_n988_ = new_n873_ & new_n959_;
  assign new_n989_ = new_n873_;
  assign new_n990_ = new_n873_;
  assign new_n991_ = new_n366_ & new_n963_;
  assign new_n992_ = new_n963_ & new_n366_;
  assign new_n993_ = ~new_n963_ & ~new_n366_;
  assign new_n994_ = ~new_n366_ & ~new_n963_;
  assign new_n995_ = new_n874_ & new_n960_;
  assign new_n996_ = new_n874_;
  assign new_n997_ = new_n874_;
  assign new_n998_ = new_n875_ & new_n961_;
  assign new_n999_ = new_n875_;
  assign new_n1000_ = new_n875_;
  assign new_n1001_ = new_n370_ & new_n964_;
  assign new_n1002_ = new_n370_ & new_n964_;
  assign new_n1003_ = new_n371_ & new_n928_;
  assign new_n1004_ = new_n371_ & new_n928_;
  assign new_n1005_ = new_n876_ & new_n923_;
  assign new_n1006_ = new_n876_;
  assign new_n1007_ = new_n876_;
  assign new_n1008_ = new_n373_ & new_n927_;
  assign new_n1009_ = new_n373_ & new_n927_;
  assign new_n1010_ = new_n877_ & new_n922_;
  assign new_n1011_ = new_n877_;
  assign new_n1012_ = new_n877_;
  assign new_n1013_ = new_n375_ & new_n926_;
  assign new_n1014_ = new_n375_ & new_n926_;
  assign new_n1015_ = new_n878_ & new_n921_;
  assign new_n1016_ = new_n878_;
  assign new_n1017_ = new_n878_;
  assign new_n1018_ = new_n377_ & new_n929_;
  assign new_n1019_ = new_n377_ & new_n929_;
  assign new_n1020_ = ~new_n377_ & ~new_n929_;
  assign new_n1021_ = new_n879_ & new_n924_;
  assign new_n1022_ = new_n879_;
  assign new_n1023_ = new_n879_;
  assign new_n1024_ = ~new_n880_;
  assign new_n1025_ = ~new_n881_;
  assign new_n1026_ = new_n882_;
  assign new_n1027_ = new_n882_;
  assign new_n1028_ = new_n883_;
  assign new_n1029_ = new_n883_;
  assign new_n1030_ = ~new_n884_;
  assign new_n1031_ = ~new_n941_ | ~new_n713_;
  assign new_n1032_ = ~new_n940_ | ~new_n715_;
  assign new_n1033_ = new_n388_ & new_n974_;
  assign new_n1034_ = new_n388_ & new_n974_;
  assign new_n1035_ = new_n885_ & new_n956_;
  assign new_n1036_ = new_n885_;
  assign new_n1037_ = new_n885_;
  assign new_n1038_ = new_n390_ & new_n967_;
  assign new_n1039_ = new_n390_ & new_n967_;
  assign new_n1040_ = new_n886_ & new_n950_;
  assign new_n1041_ = new_n886_;
  assign new_n1042_ = new_n886_;
  assign new_n1043_ = new_n392_ & new_n969_;
  assign new_n1044_ = new_n392_ & new_n969_;
  assign new_n1045_ = new_n887_ & new_n952_;
  assign new_n1046_ = new_n887_;
  assign new_n1047_ = new_n887_;
  assign new_n1048_ = new_n394_ & new_n970_;
  assign new_n1049_ = new_n394_ & new_n970_;
  assign new_n1050_ = ~new_n394_ & ~new_n970_;
  assign new_n1051_ = new_n888_ & new_n953_;
  assign new_n1052_ = new_n888_;
  assign new_n1053_ = new_n888_;
  assign new_n1054_ = ~new_n889_;
  assign new_n1055_ = ~new_n920_;
  assign new_n1056_ = new_n921_;
  assign new_n1057_ = new_n921_;
  assign new_n1058_ = new_n922_;
  assign new_n1059_ = new_n922_;
  assign new_n1060_ = new_n923_;
  assign new_n1061_ = new_n923_;
  assign new_n1062_ = new_n924_;
  assign new_n1063_ = new_n924_;
  assign new_n1064_ = ~new_n925_;
  assign new_n1065_ = new_n926_;
  assign new_n1066_ = new_n926_;
  assign new_n1067_ = new_n926_;
  assign new_n1068_ = new_n927_;
  assign new_n1069_ = new_n927_;
  assign new_n1070_ = new_n927_;
  assign new_n1071_ = new_n928_;
  assign new_n1072_ = new_n928_;
  assign new_n1073_ = new_n928_;
  assign new_n1074_ = new_n929_;
  assign new_n1075_ = new_n929_;
  assign new_n1076_ = new_n929_;
  assign new_n1077_ = new_n911_ | new_n762_;
  assign new_n1078_ = new_n895_ | new_n763_;
  assign new_n1079_ = new_n896_ | new_n764_;
  assign new_n1080_ = new_n912_ | new_n765_;
  assign new_n1081_ = new_n897_ | new_n766_;
  assign new_n1082_ = new_n913_ | new_n767_;
  assign new_n1083_ = new_n903_ | new_n768_;
  assign new_n1084_ = new_n918_ | new_n769_;
  assign new_n1085_ = new_n919_ | new_n770_;
  assign new_n1086_ = new_n909_ | new_n771_;
  assign new_n1087_ = new_n915_ | new_n772_;
  assign new_n1088_ = new_n900_ | new_n773_;
  assign new_n1089_ = new_n503_ & new_n968_;
  assign new_n1090_ = new_n503_ & new_n968_;
  assign new_n1091_ = new_n930_ & new_n951_;
  assign new_n1092_ = new_n930_;
  assign new_n1093_ = new_n930_;
  assign new_n1094_ = new_n910_ | new_n782_;
  assign new_n1095_ = new_n894_ | new_n783_;
  assign new_n1096_ = new_n898_ | new_n784_;
  assign new_n1097_ = new_n914_ | new_n785_;
  assign new_n1098_ = new_n901_ | new_n786_;
  assign new_n1099_ = new_n916_ | new_n787_;
  assign new_n1100_ = new_n902_ | new_n788_;
  assign new_n1101_ = new_n917_ | new_n789_;
  assign new_n1102_ = new_n856_ | new_n797_;
  assign new_n1103_ = new_n855_ | new_n798_;
  assign new_n1104_ = new_n854_ | new_n799_;
  assign new_n1105_ = new_n858_ | new_n800_;
  assign new_n1106_ = new_n859_ | new_n801_;
  assign new_n1107_ = new_n867_ | new_n802_;
  assign new_n1108_ = new_n866_ | new_n803_;
  assign new_n1109_ = new_n868_ | new_n804_;
  assign new_n1110_ = new_n865_ | new_n805_;
  assign new_n1111_ = new_n869_ | new_n806_;
  assign new_n1112_ = new_n870_ | new_n808_;
  assign new_n1113_ = new_n908_ | new_n809_;
  assign new_n1114_ = new_n931_;
  assign new_n1115_ = new_n931_;
  assign new_n1116_ = new_n851_ | new_n813_;
  assign new_n1117_ = new_n852_ | new_n814_;
  assign new_n1118_ = new_n853_ | new_n815_;
  assign new_n1119_ = new_n857_ | new_n816_;
  assign new_n1120_ = new_n860_ | new_n817_;
  assign new_n1121_ = new_n861_ | new_n818_;
  assign new_n1122_ = new_n862_ | new_n819_;
  assign new_n1123_ = new_n863_ | new_n820_;
  assign new_n1124_ = new_n864_ | new_n821_;
  assign new_n1125_ = new_n907_ | new_n822_;
  assign new_n1126_ = new_n932_;
  assign new_n1127_ = new_n932_;
  assign new_n1128_ = new_n933_;
  assign new_n1129_ = new_n933_;
  assign new_n1130_ = new_n904_ | new_n823_;
  assign new_n1131_ = ~new_n934_;
  assign new_n1132_ = new_n890_ | new_n824_;
  assign new_n1133_ = new_n935_;
  assign new_n1134_ = new_n899_ | new_n825_;
  assign new_n1135_ = ~new_n505_ | ~new_n850_;
  assign new_n1136_ = new_n883_ & new_n668_;
  assign new_n1137_ = new_n883_ & new_n668_;
  assign new_n1138_ = new_n883_ & new_n668_;
  assign new_n1139_ = new_n883_ & new_n668_;
  assign new_n1140_ = new_n882_ & new_n669_;
  assign new_n1141_ = new_n942_;
  assign new_n1142_ = new_n942_;
  assign new_n1143_ = new_n905_ | new_n833_;
  assign new_n1144_ = new_n906_ | new_n834_;
  assign new_n1145_ = new_n943_;
  assign new_n1146_ = new_n943_;
  assign new_n1147_ = new_n891_ | new_n835_;
  assign new_n1148_ = new_n944_;
  assign new_n1149_ = new_n944_;
  assign new_n1150_ = new_n892_ | new_n836_;
  assign new_n1151_ = new_n945_;
  assign new_n1152_ = new_n945_;
  assign new_n1153_ = new_n893_ | new_n837_;
  assign new_n1154_ = new_n946_;
  assign new_n1155_ = new_n946_;
  assign new_n1156_ = new_n947_;
  assign new_n1157_ = new_n948_;
  assign new_n1158_ = new_n948_;
  assign new_n1159_ = new_n411_ & new_n935_;
  assign new_n1160_ = ~new_n949_;
  assign new_n1161_ = new_n950_;
  assign new_n1162_ = new_n950_;
  assign new_n1163_ = new_n951_;
  assign new_n1164_ = new_n951_;
  assign new_n1165_ = new_n952_;
  assign new_n1166_ = new_n952_;
  assign new_n1167_ = new_n953_;
  assign new_n1168_ = new_n953_;
  assign new_n1169_ = ~new_n954_;
  assign new_n1170_ = ~new_n955_;
  assign new_n1171_ = new_n956_;
  assign new_n1172_ = new_n956_;
  assign new_n1173_ = new_n957_;
  assign new_n1174_ = new_n957_;
  assign new_n1175_ = new_n958_;
  assign new_n1176_ = new_n958_;
  assign new_n1177_ = new_n959_;
  assign new_n1178_ = new_n959_;
  assign new_n1179_ = new_n960_;
  assign new_n1180_ = new_n960_;
  assign new_n1181_ = new_n961_;
  assign new_n1182_ = new_n961_;
  assign new_n1183_ = new_n962_;
  assign new_n1184_ = new_n962_;
  assign new_n1185_ = new_n962_;
  assign new_n1186_ = new_n963_;
  assign new_n1187_ = new_n963_;
  assign new_n1188_ = new_n963_;
  assign new_n1189_ = new_n964_;
  assign new_n1190_ = new_n964_;
  assign new_n1191_ = new_n964_;
  assign new_n1192_ = new_n965_;
  assign new_n1193_ = new_n965_;
  assign new_n1194_ = new_n965_;
  assign new_n1195_ = new_n966_;
  assign new_n1196_ = new_n966_;
  assign new_n1197_ = new_n966_;
  assign new_n1198_ = new_n967_;
  assign new_n1199_ = new_n967_;
  assign new_n1200_ = new_n967_;
  assign new_n1201_ = new_n968_;
  assign new_n1202_ = new_n968_;
  assign new_n1203_ = new_n968_;
  assign new_n1204_ = new_n969_;
  assign new_n1205_ = new_n969_;
  assign new_n1206_ = new_n969_;
  assign new_n1207_ = new_n970_;
  assign new_n1208_ = new_n970_;
  assign new_n1209_ = new_n970_;
  assign new_n1210_ = ~new_n971_;
  assign new_n1211_ = ~new_n972_;
  assign new_n1212_ = ~new_n973_;
  assign new_n1213_ = new_n974_;
  assign new_n1214_ = new_n974_;
  assign new_n1215_ = new_n974_;
  assign new_n1216_ = new_n318_ & new_n1113_;
  assign new_n1217_ = new_n318_ & new_n1113_;
  assign new_n1218_ = new_n320_ & new_n1125_;
  assign new_n1219_ = new_n320_ & new_n1125_;
  assign new_n1220_ = new_n322_ & new_n1144_;
  assign new_n1221_ = new_n322_ & new_n1144_;
  assign new_n1222_ = new_n1143_ & new_n324_;
  assign new_n1223_ = new_n324_ & new_n1143_;
  assign new_n1224_ = ~new_n324_ & ~new_n1143_;
  assign new_n1225_ = ~new_n1143_ & ~new_n324_;
  assign new_n1226_ = new_n326_ & new_n1130_;
  assign new_n1227_ = new_n326_ & new_n1130_;
  assign new_n1228_ = new_n328_ & new_n1083_;
  assign new_n1229_ = new_n328_ & new_n1083_;
  assign new_n1230_ = new_n330_ & new_n1100_;
  assign new_n1231_ = new_n330_ & new_n1100_;
  assign new_n1232_ = new_n332_ & new_n1098_;
  assign new_n1233_ = new_n332_ & new_n1098_;
  assign new_n1234_ = new_n334_ & new_n1086_;
  assign new_n1235_ = new_n334_ & new_n1086_;
  assign new_n1236_ = ~new_n334_ & ~new_n1086_;
  assign new_n1237_ = new_n338_ & new_n1096_;
  assign new_n1238_ = new_n338_ & new_n1096_;
  assign new_n1239_ = new_n340_ & new_n1081_;
  assign new_n1240_ = new_n340_ & new_n1081_;
  assign new_n1241_ = new_n342_ & new_n1079_;
  assign new_n1242_ = new_n342_ & new_n1079_;
  assign new_n1243_ = new_n1078_ & new_n344_;
  assign new_n1244_ = new_n344_ & new_n1078_;
  assign new_n1245_ = ~new_n344_ & ~new_n1078_;
  assign new_n1246_ = ~new_n1078_ & ~new_n344_;
  assign new_n1247_ = new_n346_ & new_n1095_;
  assign new_n1248_ = new_n346_ & new_n1095_;
  assign new_n1249_ = new_n348_ & new_n1153_;
  assign new_n1250_ = new_n348_ & new_n1153_;
  assign new_n1251_ = new_n350_ & new_n1150_;
  assign new_n1252_ = new_n350_ & new_n1150_;
  assign new_n1253_ = new_n352_ & new_n1147_;
  assign new_n1254_ = new_n352_ & new_n1147_;
  assign new_n1255_ = ~new_n977_;
  assign new_n1256_ = ~new_n978_;
  assign new_n1257_ = ~new_n1193_ | ~new_n575_;
  assign new_n1258_ = ~new_n1194_ | ~new_n576_;
  assign new_n1259_ = ~new_n982_;
  assign new_n1260_ = ~new_n983_;
  assign new_n1261_ = ~new_n1195_ | ~new_n578_;
  assign new_n1262_ = ~new_n1196_ | ~new_n579_;
  assign new_n1263_ = ~new_n989_;
  assign new_n1264_ = ~new_n990_;
  assign new_n1265_ = ~new_n1185_ | ~new_n581_;
  assign new_n1266_ = ~new_n1184_ | ~new_n582_;
  assign new_n1267_ = new_n991_;
  assign new_n1268_ = new_n992_;
  assign new_n1269_ = ~new_n1187_ | ~new_n583_;
  assign new_n1270_ = ~new_n993_;
  assign new_n1271_ = ~new_n994_;
  assign new_n1272_ = ~new_n1186_ | ~new_n584_;
  assign new_n1273_ = ~new_n996_;
  assign new_n1274_ = ~new_n997_;
  assign new_n1275_ = ~new_n999_;
  assign new_n1276_ = ~new_n1000_;
  assign new_n1277_ = ~new_n1191_ | ~new_n587_;
  assign new_n1278_ = ~new_n1190_ | ~new_n588_;
  assign new_n1279_ = ~new_n1073_ | ~new_n589_;
  assign new_n1280_ = ~new_n1072_ | ~new_n590_;
  assign new_n1281_ = ~new_n1006_;
  assign new_n1282_ = ~new_n1007_;
  assign new_n1283_ = ~new_n1011_;
  assign new_n1284_ = ~new_n1012_;
  assign new_n1285_ = ~new_n1070_ | ~new_n593_;
  assign new_n1286_ = ~new_n1069_ | ~new_n594_;
  assign new_n1287_ = ~new_n1067_ | ~new_n595_;
  assign new_n1288_ = ~new_n1066_ | ~new_n596_;
  assign new_n1289_ = ~new_n1016_;
  assign new_n1290_ = ~new_n1017_;
  assign new_n1291_ = new_n1018_;
  assign new_n1292_ = ~new_n1020_;
  assign new_n1293_ = ~new_n1076_ | ~new_n598_;
  assign new_n1294_ = ~new_n1022_ | ~new_n1024_;
  assign new_n1295_ = ~new_n1022_;
  assign new_n1296_ = ~new_n1023_;
  assign new_n1297_ = ~new_n1075_ | ~new_n600_;
  assign new_n1298_ = ~new_n881_ | ~new_n1030_;
  assign new_n1299_ = new_n479_ | new_n1139_;
  assign new_n1300_ = ~new_n479_ & ~new_n1138_;
  assign new_n1301_ = new_n479_ | new_n1137_;
  assign new_n1302_ = new_n480_ | new_n1140_;
  assign new_n1303_ = ~new_n1026_;
  assign new_n1304_ = ~new_n1027_;
  assign new_n1305_ = new_n1032_ & new_n882_;
  assign new_n1306_ = new_n1031_ & new_n883_;
  assign new_n1307_ = ~new_n1028_;
  assign new_n1308_ = new_n1031_ & new_n883_;
  assign new_n1309_ = new_n1031_ & new_n883_;
  assign new_n1310_ = ~new_n1029_;
  assign new_n1311_ = ~new_n884_ | ~new_n1025_;
  assign new_n1312_ = new_n1031_;
  assign new_n1313_ = new_n1031_;
  assign new_n1314_ = ~new_n1032_;
  assign new_n1315_ = ~new_n1036_;
  assign new_n1316_ = ~new_n1037_;
  assign new_n1317_ = ~new_n1214_ | ~new_n609_;
  assign new_n1318_ = ~new_n1215_ | ~new_n610_;
  assign new_n1319_ = ~new_n1198_ | ~new_n611_;
  assign new_n1320_ = ~new_n1199_ | ~new_n612_;
  assign new_n1321_ = ~new_n1041_;
  assign new_n1322_ = ~new_n1042_;
  assign new_n1323_ = ~new_n1204_ | ~new_n614_;
  assign new_n1324_ = ~new_n1046_;
  assign new_n1325_ = ~new_n1047_;
  assign new_n1326_ = ~new_n1205_ | ~new_n616_;
  assign new_n1327_ = new_n1048_;
  assign new_n1328_ = ~new_n1050_;
  assign new_n1329_ = ~new_n1208_ | ~new_n617_;
  assign new_n1330_ = ~new_n1052_ | ~new_n1054_;
  assign new_n1331_ = ~new_n1052_;
  assign new_n1332_ = ~new_n1053_;
  assign new_n1333_ = ~new_n1209_ | ~new_n619_;
  assign new_n1334_ = ~new_n1062_ | ~new_n1055_;
  assign new_n1335_ = ~new_n1056_;
  assign new_n1336_ = ~new_n1057_;
  assign new_n1337_ = ~new_n1058_;
  assign new_n1338_ = ~new_n1059_;
  assign new_n1339_ = ~new_n1060_;
  assign new_n1340_ = ~new_n1061_;
  assign new_n1341_ = ~new_n1062_;
  assign new_n1342_ = ~new_n1063_;
  assign new_n1343_ = ~new_n1074_ | ~new_n1064_;
  assign new_n1344_ = ~new_n1065_;
  assign new_n1345_ = ~new_n1066_;
  assign new_n1346_ = ~new_n1067_;
  assign new_n1347_ = ~new_n1068_;
  assign new_n1348_ = ~new_n1069_;
  assign new_n1349_ = ~new_n1070_;
  assign new_n1350_ = ~new_n1071_;
  assign new_n1351_ = ~new_n1072_;
  assign new_n1352_ = ~new_n1073_;
  assign new_n1353_ = ~new_n1074_;
  assign new_n1354_ = ~new_n1075_;
  assign new_n1355_ = ~new_n1076_;
  assign new_n1356_ = new_n1077_;
  assign new_n1357_ = new_n1124_ & new_n1077_;
  assign new_n1358_ = new_n1077_;
  assign new_n1359_ = new_n1078_;
  assign new_n1360_ = new_n1078_;
  assign new_n1361_ = new_n1078_;
  assign new_n1362_ = new_n1079_;
  assign new_n1363_ = new_n1079_;
  assign new_n1364_ = new_n1079_;
  assign new_n1365_ = new_n1123_ & new_n1080_;
  assign new_n1366_ = new_n1080_;
  assign new_n1367_ = new_n1080_;
  assign new_n1368_ = new_n1081_;
  assign new_n1369_ = new_n1081_;
  assign new_n1370_ = new_n1081_;
  assign new_n1371_ = new_n1122_ & new_n1082_;
  assign new_n1372_ = new_n1082_;
  assign new_n1373_ = new_n1082_;
  assign new_n1374_ = new_n1083_;
  assign new_n1375_ = new_n1083_;
  assign new_n1376_ = new_n1083_;
  assign new_n1377_ = new_n1102_ & new_n1084_;
  assign new_n1378_ = new_n1084_;
  assign new_n1379_ = new_n1084_;
  assign new_n1380_ = new_n1106_ & new_n1085_;
  assign new_n1381_ = new_n1085_;
  assign new_n1382_ = new_n1085_;
  assign new_n1383_ = new_n1086_;
  assign new_n1384_ = new_n1086_;
  assign new_n1385_ = new_n1086_;
  assign new_n1386_ = ~new_n1087_;
  assign new_n1387_ = ~new_n1088_;
  assign new_n1388_ = ~new_n1202_ | ~new_n780_;
  assign new_n1389_ = ~new_n1203_ | ~new_n781_;
  assign new_n1390_ = ~new_n1092_;
  assign new_n1391_ = ~new_n1093_;
  assign new_n1392_ = new_n1094_;
  assign new_n1393_ = new_n1110_ & new_n1094_;
  assign new_n1394_ = new_n1094_;
  assign new_n1395_ = new_n1095_;
  assign new_n1396_ = new_n1095_;
  assign new_n1397_ = new_n1095_;
  assign new_n1398_ = new_n1096_;
  assign new_n1399_ = new_n1096_;
  assign new_n1400_ = new_n1096_;
  assign new_n1401_ = new_n1097_;
  assign new_n1402_ = new_n1121_ & new_n1097_;
  assign new_n1403_ = new_n1097_;
  assign new_n1404_ = new_n1098_;
  assign new_n1405_ = new_n1098_;
  assign new_n1406_ = new_n1098_;
  assign new_n1407_ = new_n1105_ & new_n1099_;
  assign new_n1408_ = new_n1099_;
  assign new_n1409_ = new_n1099_;
  assign new_n1410_ = new_n1100_;
  assign new_n1411_ = new_n1100_;
  assign new_n1412_ = new_n1100_;
  assign new_n1413_ = new_n1101_;
  assign new_n1414_ = new_n1119_ & new_n1101_;
  assign new_n1415_ = new_n1101_;
  assign new_n1416_ = new_n1102_;
  assign new_n1417_ = new_n1102_;
  assign new_n1418_ = new_n1103_;
  assign new_n1419_ = new_n1103_;
  assign new_n1420_ = new_n1104_;
  assign new_n1421_ = new_n1104_;
  assign new_n1422_ = new_n1105_;
  assign new_n1423_ = new_n1105_;
  assign new_n1424_ = new_n1106_;
  assign new_n1425_ = new_n1106_;
  assign new_n1426_ = new_n1107_;
  assign new_n1427_ = new_n1107_;
  assign new_n1428_ = new_n1108_;
  assign new_n1429_ = new_n1108_;
  assign new_n1430_ = new_n1109_;
  assign new_n1431_ = new_n1109_;
  assign new_n1432_ = new_n1110_;
  assign new_n1433_ = new_n1110_;
  assign new_n1434_ = ~new_n1111_;
  assign new_n1435_ = ~new_n1112_;
  assign new_n1436_ = new_n1113_;
  assign new_n1437_ = new_n1113_;
  assign new_n1438_ = new_n1113_;
  assign new_n1439_ = new_n1116_ & new_n931_;
  assign new_n1440_ = ~new_n1114_;
  assign new_n1441_ = ~new_n1115_;
  assign new_n1442_ = new_n1116_;
  assign new_n1443_ = new_n1116_;
  assign new_n1444_ = new_n1117_;
  assign new_n1445_ = new_n1117_;
  assign new_n1446_ = new_n1118_;
  assign new_n1447_ = new_n1118_;
  assign new_n1448_ = new_n1119_;
  assign new_n1449_ = new_n1119_;
  assign new_n1450_ = ~new_n1120_;
  assign new_n1451_ = new_n1121_;
  assign new_n1452_ = new_n1121_;
  assign new_n1453_ = new_n1122_;
  assign new_n1454_ = new_n1122_;
  assign new_n1455_ = new_n1123_;
  assign new_n1456_ = new_n1123_;
  assign new_n1457_ = new_n1124_;
  assign new_n1458_ = new_n1124_;
  assign new_n1459_ = new_n1125_;
  assign new_n1460_ = new_n1125_;
  assign new_n1461_ = new_n1125_;
  assign new_n1462_ = new_n1117_ & new_n932_;
  assign new_n1463_ = ~new_n1126_;
  assign new_n1464_ = ~new_n1127_;
  assign new_n1465_ = new_n1103_ & new_n933_;
  assign new_n1466_ = ~new_n1128_;
  assign new_n1467_ = ~new_n1129_;
  assign new_n1468_ = new_n1130_;
  assign new_n1469_ = new_n1130_;
  assign new_n1470_ = new_n1130_;
  assign new_n1471_ = ~new_n1133_ | ~new_n1131_;
  assign new_n1472_ = ~new_n1132_;
  assign new_n1473_ = ~new_n1133_;
  assign new_n1474_ = new_n1134_;
  assign new_n1475_ = new_n975_ & new_n826_;
  assign new_n1476_ = ~new_n1135_ | ~new_n936_;
  assign new_n1477_ = ~new_n1026_ | ~new_n939_;
  assign new_n1478_ = ~new_n1027_ | ~new_n829_;
  assign new_n1479_ = new_n1104_ & new_n942_;
  assign new_n1480_ = ~new_n1141_;
  assign new_n1481_ = ~new_n1142_;
  assign new_n1482_ = new_n1143_;
  assign new_n1483_ = new_n1143_;
  assign new_n1484_ = new_n1143_;
  assign new_n1485_ = new_n1144_;
  assign new_n1486_ = new_n1144_;
  assign new_n1487_ = new_n1144_;
  assign new_n1488_ = new_n1118_ & new_n943_;
  assign new_n1489_ = ~new_n1145_;
  assign new_n1490_ = ~new_n1146_;
  assign new_n1491_ = new_n1147_;
  assign new_n1492_ = new_n1147_;
  assign new_n1493_ = new_n1147_;
  assign new_n1494_ = new_n1109_ & new_n944_;
  assign new_n1495_ = ~new_n1148_;
  assign new_n1496_ = ~new_n1149_;
  assign new_n1497_ = new_n1150_;
  assign new_n1498_ = new_n1150_;
  assign new_n1499_ = new_n1150_;
  assign new_n1500_ = ~new_n1151_;
  assign new_n1501_ = new_n1107_ & new_n945_;
  assign new_n1502_ = ~new_n1152_;
  assign new_n1503_ = new_n1153_;
  assign new_n1504_ = new_n1153_;
  assign new_n1505_ = new_n1153_;
  assign new_n1506_ = new_n1108_ & new_n946_;
  assign new_n1507_ = ~new_n1154_;
  assign new_n1508_ = ~new_n1155_;
  assign new_n1509_ = new_n947_ & new_n1159_;
  assign new_n1510_ = ~new_n1156_;
  assign new_n1511_ = ~new_n1157_;
  assign new_n1512_ = ~new_n1158_;
  assign new_n1513_ = new_n1159_;
  assign new_n1514_ = new_n1134_ & new_n411_;
  assign new_n1515_ = ~new_n1160_;
  assign new_n1516_ = ~new_n1161_;
  assign new_n1517_ = ~new_n1162_;
  assign new_n1518_ = ~new_n1163_;
  assign new_n1519_ = ~new_n1164_;
  assign new_n1520_ = ~new_n1165_;
  assign new_n1521_ = ~new_n1166_;
  assign new_n1522_ = ~new_n1167_;
  assign new_n1523_ = ~new_n1168_;
  assign new_n1524_ = ~new_n954_ | ~new_n1170_;
  assign new_n1525_ = ~new_n955_ | ~new_n1169_;
  assign new_n1526_ = ~new_n1171_;
  assign new_n1527_ = ~new_n1172_;
  assign new_n1528_ = ~new_n1173_;
  assign new_n1529_ = ~new_n1174_;
  assign new_n1530_ = ~new_n1175_;
  assign new_n1531_ = ~new_n1176_;
  assign new_n1532_ = ~new_n1177_;
  assign new_n1533_ = ~new_n1178_;
  assign new_n1534_ = ~new_n1179_;
  assign new_n1535_ = ~new_n1180_;
  assign new_n1536_ = ~new_n1181_;
  assign new_n1537_ = ~new_n1182_;
  assign new_n1538_ = ~new_n1183_;
  assign new_n1539_ = ~new_n1184_;
  assign new_n1540_ = ~new_n1185_;
  assign new_n1541_ = ~new_n1186_;
  assign new_n1542_ = ~new_n1187_;
  assign new_n1543_ = ~new_n1188_;
  assign new_n1544_ = ~new_n1189_;
  assign new_n1545_ = ~new_n1190_;
  assign new_n1546_ = ~new_n1191_;
  assign new_n1547_ = ~new_n1192_;
  assign new_n1548_ = ~new_n1193_;
  assign new_n1549_ = ~new_n1194_;
  assign new_n1550_ = ~new_n1195_;
  assign new_n1551_ = ~new_n1196_;
  assign new_n1552_ = ~new_n1197_;
  assign new_n1553_ = ~new_n1198_;
  assign new_n1554_ = ~new_n1199_;
  assign new_n1555_ = ~new_n1200_;
  assign new_n1556_ = ~new_n1201_;
  assign new_n1557_ = ~new_n1202_;
  assign new_n1558_ = ~new_n1203_;
  assign new_n1559_ = ~new_n1204_;
  assign new_n1560_ = ~new_n1205_;
  assign new_n1561_ = ~new_n1206_;
  assign new_n1562_ = ~new_n1207_;
  assign new_n1563_ = ~new_n1208_;
  assign new_n1564_ = ~new_n1209_;
  assign new_n1565_ = ~new_n1210_;
  assign new_n1566_ = ~new_n972_ | ~new_n1212_;
  assign new_n1567_ = ~new_n973_ | ~new_n1211_;
  assign new_n1568_ = ~new_n1213_;
  assign new_n1569_ = ~new_n1214_;
  assign new_n1570_ = ~new_n1215_;
  assign new_n1571_ = new_n1476_ & new_n975_;
  assign new_n1572_ = ~new_n1436_ | ~new_n540_;
  assign new_n1573_ = ~new_n1438_ | ~new_n541_;
  assign new_n1574_ = ~new_n1459_ | ~new_n542_;
  assign new_n1575_ = ~new_n1461_ | ~new_n543_;
  assign new_n1576_ = ~new_n1487_ | ~new_n544_;
  assign new_n1577_ = ~new_n1486_ | ~new_n545_;
  assign new_n1578_ = new_n1222_;
  assign new_n1579_ = new_n1223_;
  assign new_n1580_ = ~new_n1224_;
  assign new_n1581_ = ~new_n1483_ | ~new_n546_;
  assign new_n1582_ = ~new_n1484_ | ~new_n547_;
  assign new_n1583_ = ~new_n1225_;
  assign new_n1584_ = ~new_n1470_ | ~new_n548_;
  assign new_n1585_ = ~new_n1468_ | ~new_n549_;
  assign new_n1586_ = ~new_n1375_ | ~new_n550_;
  assign new_n1587_ = ~new_n1376_ | ~new_n551_;
  assign new_n1588_ = ~new_n1411_ | ~new_n552_;
  assign new_n1589_ = ~new_n1412_ | ~new_n553_;
  assign new_n1590_ = ~new_n1405_ | ~new_n554_;
  assign new_n1591_ = ~new_n1406_ | ~new_n555_;
  assign new_n1592_ = new_n1235_;
  assign new_n1593_ = ~new_n1384_ | ~new_n556_;
  assign new_n1594_ = ~new_n1236_;
  assign new_n1595_ = ~new_n1385_ | ~new_n557_;
  assign new_n1596_ = ~new_n1399_ | ~new_n558_;
  assign new_n1597_ = ~new_n1400_ | ~new_n559_;
  assign new_n1598_ = ~new_n1368_ | ~new_n560_;
  assign new_n1599_ = ~new_n1369_ | ~new_n561_;
  assign new_n1600_ = ~new_n1363_ | ~new_n562_;
  assign new_n1601_ = ~new_n1364_ | ~new_n563_;
  assign new_n1602_ = new_n1243_;
  assign new_n1603_ = new_n1244_;
  assign new_n1604_ = ~new_n1245_;
  assign new_n1605_ = ~new_n1360_ | ~new_n564_;
  assign new_n1606_ = ~new_n1359_ | ~new_n565_;
  assign new_n1607_ = ~new_n1246_;
  assign new_n1608_ = ~new_n1397_ | ~new_n566_;
  assign new_n1609_ = ~new_n1396_ | ~new_n567_;
  assign new_n1610_ = ~new_n1504_ | ~new_n568_;
  assign new_n1611_ = ~new_n1503_ | ~new_n569_;
  assign new_n1612_ = ~new_n1499_ | ~new_n570_;
  assign new_n1613_ = ~new_n1498_ | ~new_n571_;
  assign new_n1614_ = ~new_n1492_ | ~new_n572_;
  assign new_n1615_ = ~new_n1491_ | ~new_n573_;
  assign new_n1616_ = ~new_n977_ | ~new_n1259_;
  assign new_n1617_ = ~new_n978_ | ~new_n1529_;
  assign new_n1618_ = ~new_n461_ | ~new_n1548_;
  assign new_n1619_ = ~new_n462_ | ~new_n1549_;
  assign new_n1620_ = ~new_n982_ | ~new_n1255_;
  assign new_n1621_ = ~new_n983_ | ~new_n1530_;
  assign new_n1622_ = ~new_n463_ | ~new_n1550_;
  assign new_n1623_ = ~new_n464_ | ~new_n1551_;
  assign new_n1624_ = ~new_n989_ | ~new_n1533_;
  assign new_n1625_ = ~new_n990_ | ~new_n1273_;
  assign new_n1626_ = ~new_n465_ | ~new_n1540_;
  assign new_n1627_ = ~new_n466_ | ~new_n1539_;
  assign new_n1628_ = ~new_n1267_;
  assign new_n1629_ = ~new_n1268_;
  assign new_n1630_ = ~new_n467_ | ~new_n1542_;
  assign new_n1631_ = ~new_n468_ | ~new_n1541_;
  assign new_n1632_ = ~new_n996_ | ~new_n1264_;
  assign new_n1633_ = ~new_n997_ | ~new_n1534_;
  assign new_n1634_ = ~new_n999_ | ~new_n1282_;
  assign new_n1635_ = ~new_n1000_ | ~new_n1537_;
  assign new_n1636_ = ~new_n469_ | ~new_n1546_;
  assign new_n1637_ = ~new_n470_ | ~new_n1545_;
  assign new_n1638_ = ~new_n471_ | ~new_n1352_;
  assign new_n1639_ = ~new_n472_ | ~new_n1351_;
  assign new_n1640_ = ~new_n1006_ | ~new_n1339_;
  assign new_n1641_ = ~new_n1007_ | ~new_n1275_;
  assign new_n1642_ = ~new_n1011_ | ~new_n1290_;
  assign new_n1643_ = ~new_n1012_ | ~new_n1338_;
  assign new_n1644_ = ~new_n473_ | ~new_n1349_;
  assign new_n1645_ = ~new_n474_ | ~new_n1348_;
  assign new_n1646_ = ~new_n475_ | ~new_n1346_;
  assign new_n1647_ = ~new_n476_ | ~new_n1345_;
  assign new_n1648_ = ~new_n1016_ | ~new_n1335_;
  assign new_n1649_ = ~new_n1017_ | ~new_n1283_;
  assign new_n1650_ = ~new_n1291_;
  assign new_n1651_ = ~new_n477_ | ~new_n1355_;
  assign new_n1652_ = ~new_n1023_ | ~new_n1342_;
  assign new_n1653_ = ~new_n478_ | ~new_n1354_;
  assign new_n1654_ = ~new_n880_ | ~new_n1295_;
  assign new_n1655_ = ~new_n1311_ | ~new_n1298_;
  assign new_n1656_ = new_n1299_ | new_n1306_;
  assign new_n1657_ = ~new_n1299_;
  assign new_n1658_ = ~new_n1300_;
  assign new_n1659_ = ~new_n1301_;
  assign new_n1660_ = new_n1309_ | new_n479_ | new_n1136_;
  assign new_n1661_ = ~new_n1302_;
  assign new_n1662_ = ~new_n1305_;
  assign new_n1663_ = ~new_n1308_;
  assign new_n1664_ = ~new_n1312_;
  assign new_n1665_ = ~new_n1313_;
  assign new_n1666_ = ~new_n1036_ | ~new_n1322_;
  assign new_n1667_ = ~new_n1037_ | ~new_n1527_;
  assign new_n1668_ = ~new_n484_ | ~new_n1569_;
  assign new_n1669_ = ~new_n485_ | ~new_n1570_;
  assign new_n1670_ = ~new_n486_ | ~new_n1553_;
  assign new_n1671_ = ~new_n487_ | ~new_n1554_;
  assign new_n1672_ = ~new_n1041_ | ~new_n1517_;
  assign new_n1673_ = ~new_n1042_ | ~new_n1315_;
  assign new_n1674_ = ~new_n488_ | ~new_n1559_;
  assign new_n1675_ = ~new_n1046_ | ~new_n1521_;
  assign new_n1676_ = ~new_n1047_ | ~new_n1390_;
  assign new_n1677_ = ~new_n489_ | ~new_n1560_;
  assign new_n1678_ = ~new_n1327_;
  assign new_n1679_ = ~new_n490_ | ~new_n1563_;
  assign new_n1680_ = ~new_n1053_ | ~new_n1523_;
  assign new_n1681_ = ~new_n491_ | ~new_n1564_;
  assign new_n1682_ = ~new_n889_ | ~new_n1331_;
  assign new_n1683_ = ~new_n920_ | ~new_n1341_;
  assign new_n1684_ = ~new_n1056_ | ~new_n1289_;
  assign new_n1685_ = ~new_n1057_ | ~new_n1337_;
  assign new_n1686_ = ~new_n1058_ | ~new_n1336_;
  assign new_n1687_ = ~new_n1059_ | ~new_n1284_;
  assign new_n1688_ = ~new_n1060_ | ~new_n1281_;
  assign new_n1689_ = ~new_n1061_ | ~new_n1536_;
  assign new_n1690_ = ~new_n1063_ | ~new_n1296_;
  assign new_n1691_ = ~new_n925_ | ~new_n1353_;
  assign new_n1692_ = ~new_n1065_ | ~new_n1347_;
  assign new_n1693_ = ~new_n1068_ | ~new_n1344_;
  assign new_n1694_ = ~new_n1071_ | ~new_n1544_;
  assign new_n1695_ = ~new_n1356_;
  assign new_n1696_ = ~new_n1358_;
  assign new_n1697_ = ~new_n1359_;
  assign new_n1698_ = ~new_n1360_;
  assign new_n1699_ = ~new_n1361_;
  assign new_n1700_ = ~new_n1362_;
  assign new_n1701_ = ~new_n1363_;
  assign new_n1702_ = ~new_n1364_;
  assign new_n1703_ = ~new_n1366_;
  assign new_n1704_ = ~new_n1367_;
  assign new_n1705_ = ~new_n1368_;
  assign new_n1706_ = ~new_n1369_;
  assign new_n1707_ = ~new_n1370_;
  assign new_n1708_ = ~new_n1372_;
  assign new_n1709_ = ~new_n1373_;
  assign new_n1710_ = ~new_n1374_;
  assign new_n1711_ = ~new_n1375_;
  assign new_n1712_ = ~new_n1376_;
  assign new_n1713_ = ~new_n1378_;
  assign new_n1714_ = ~new_n1379_ | ~new_n1467_;
  assign new_n1715_ = ~new_n1379_;
  assign new_n1716_ = ~new_n1381_;
  assign new_n1717_ = ~new_n1382_ | ~new_n1386_;
  assign new_n1718_ = ~new_n1382_;
  assign new_n1719_ = ~new_n1383_ | ~new_n1387_;
  assign new_n1720_ = ~new_n1383_;
  assign new_n1721_ = ~new_n1384_;
  assign new_n1722_ = ~new_n1385_;
  assign new_n1723_ = ~new_n657_ | ~new_n1557_;
  assign new_n1724_ = ~new_n658_ | ~new_n1558_;
  assign new_n1725_ = ~new_n1092_ | ~new_n1325_;
  assign new_n1726_ = ~new_n1093_ | ~new_n1519_;
  assign new_n1727_ = ~new_n1392_;
  assign new_n1728_ = ~new_n1394_ | ~new_n1508_;
  assign new_n1729_ = ~new_n1394_;
  assign new_n1730_ = ~new_n1395_;
  assign new_n1731_ = ~new_n1396_;
  assign new_n1732_ = ~new_n1397_;
  assign new_n1733_ = ~new_n1398_;
  assign new_n1734_ = ~new_n1399_;
  assign new_n1735_ = ~new_n1400_;
  assign new_n1736_ = ~new_n1401_;
  assign new_n1737_ = ~new_n1403_;
  assign new_n1738_ = ~new_n1404_;
  assign new_n1739_ = ~new_n1405_;
  assign new_n1740_ = ~new_n1406_;
  assign new_n1741_ = ~new_n1408_;
  assign new_n1742_ = ~new_n1409_;
  assign new_n1743_ = ~new_n1410_;
  assign new_n1744_ = ~new_n1411_;
  assign new_n1745_ = ~new_n1412_;
  assign new_n1746_ = ~new_n1413_;
  assign new_n1747_ = ~new_n1415_;
  assign new_n1748_ = ~new_n1416_;
  assign new_n1749_ = ~new_n1417_;
  assign new_n1750_ = ~new_n1418_ | ~new_n1466_;
  assign new_n1751_ = ~new_n1418_;
  assign new_n1752_ = ~new_n1419_;
  assign new_n1753_ = ~new_n1420_ | ~new_n1480_;
  assign new_n1754_ = ~new_n1420_;
  assign new_n1755_ = ~new_n1421_;
  assign new_n1756_ = ~new_n1422_;
  assign new_n1757_ = ~new_n1423_;
  assign new_n1758_ = ~new_n1424_;
  assign new_n1759_ = ~new_n1425_ | ~new_n1450_;
  assign new_n1760_ = ~new_n1425_;
  assign new_n1761_ = ~new_n1426_;
  assign new_n1762_ = ~new_n1427_ | ~new_n1500_;
  assign new_n1763_ = ~new_n1427_;
  assign new_n1764_ = ~new_n1428_ | ~new_n1507_;
  assign new_n1765_ = ~new_n1428_;
  assign new_n1766_ = ~new_n1429_;
  assign new_n1767_ = ~new_n1430_ | ~new_n1495_;
  assign new_n1768_ = ~new_n1430_;
  assign new_n1769_ = ~new_n1431_;
  assign new_n1770_ = ~new_n1432_;
  assign new_n1771_ = ~new_n1433_;
  assign new_n1772_ = ~new_n1111_ | ~new_n1435_;
  assign new_n1773_ = ~new_n1112_ | ~new_n1434_;
  assign new_n1774_ = ~new_n1436_;
  assign new_n1775_ = ~new_n1437_;
  assign new_n1776_ = ~new_n1438_;
  assign new_n1777_ = ~new_n1114_ | ~new_n1464_;
  assign new_n1778_ = ~new_n1442_ | ~new_n1441_;
  assign new_n1779_ = ~new_n1442_;
  assign new_n1780_ = ~new_n1443_;
  assign new_n1781_ = ~new_n1444_ | ~new_n1463_;
  assign new_n1782_ = ~new_n1444_;
  assign new_n1783_ = ~new_n1445_;
  assign new_n1784_ = ~new_n1446_ | ~new_n1489_;
  assign new_n1785_ = ~new_n1446_;
  assign new_n1786_ = ~new_n1447_;
  assign new_n1787_ = ~new_n1448_;
  assign new_n1788_ = ~new_n1449_;
  assign new_n1789_ = ~new_n1451_;
  assign new_n1790_ = ~new_n1452_;
  assign new_n1791_ = ~new_n1453_;
  assign new_n1792_ = ~new_n1454_;
  assign new_n1793_ = ~new_n1455_;
  assign new_n1794_ = ~new_n1456_;
  assign new_n1795_ = ~new_n1457_;
  assign new_n1796_ = ~new_n1458_;
  assign new_n1797_ = ~new_n1459_;
  assign new_n1798_ = ~new_n1460_;
  assign new_n1799_ = ~new_n1461_;
  assign new_n1800_ = ~new_n1127_ | ~new_n1440_;
  assign new_n1801_ = ~new_n1468_;
  assign new_n1802_ = ~new_n1469_;
  assign new_n1803_ = ~new_n1470_;
  assign new_n1804_ = ~new_n934_ | ~new_n1473_;
  assign new_n1805_ = ~new_n1474_ | ~new_n1472_;
  assign new_n1806_ = ~new_n1474_;
  assign new_n1807_ = new_n666_ | new_n1475_;
  assign new_n1808_ = ~new_n828_ | ~new_n1303_;
  assign new_n1809_ = ~new_n670_ | ~new_n1304_;
  assign new_n1810_ = ~new_n1142_ | ~new_n1490_;
  assign new_n1811_ = ~new_n1482_;
  assign new_n1812_ = ~new_n1483_;
  assign new_n1813_ = ~new_n1484_;
  assign new_n1814_ = ~new_n1485_;
  assign new_n1815_ = ~new_n1486_;
  assign new_n1816_ = ~new_n1487_;
  assign new_n1817_ = ~new_n1146_ | ~new_n1481_;
  assign new_n1818_ = ~new_n1491_;
  assign new_n1819_ = ~new_n1492_;
  assign new_n1820_ = ~new_n1493_;
  assign new_n1821_ = ~new_n1149_ | ~new_n1502_;
  assign new_n1822_ = ~new_n1497_;
  assign new_n1823_ = ~new_n1498_;
  assign new_n1824_ = ~new_n1499_;
  assign new_n1825_ = ~new_n1152_ | ~new_n1496_;
  assign new_n1826_ = ~new_n1503_;
  assign new_n1827_ = ~new_n1504_;
  assign new_n1828_ = ~new_n1505_;
  assign new_n1829_ = ~new_n1513_ | ~new_n1510_;
  assign new_n1830_ = new_n948_ & new_n1514_;
  assign new_n1831_ = new_n948_ & new_n1514_;
  assign new_n1832_ = ~new_n948_ & ~new_n1514_;
  assign new_n1833_ = ~new_n1513_;
  assign new_n1834_ = new_n1514_;
  assign new_n1835_ = new_n1514_;
  assign new_n1836_ = ~new_n1160_ | ~new_n1522_;
  assign new_n1837_ = ~new_n1161_ | ~new_n1526_;
  assign new_n1838_ = ~new_n1162_ | ~new_n1321_;
  assign new_n1839_ = ~new_n1163_ | ~new_n1520_;
  assign new_n1840_ = ~new_n1164_ | ~new_n1391_;
  assign new_n1841_ = ~new_n1165_ | ~new_n1518_;
  assign new_n1842_ = ~new_n1166_ | ~new_n1324_;
  assign new_n1843_ = ~new_n1167_ | ~new_n1515_;
  assign new_n1844_ = ~new_n1168_ | ~new_n1332_;
  assign new_n1845_ = ~new_n1525_ | ~new_n1524_;
  assign new_n1846_ = ~new_n1171_ | ~new_n1516_;
  assign new_n1847_ = ~new_n1172_ | ~new_n1316_;
  assign new_n1848_ = ~new_n1173_ | ~new_n1531_;
  assign new_n1849_ = ~new_n1174_ | ~new_n1256_;
  assign new_n1850_ = ~new_n1175_ | ~new_n1260_;
  assign new_n1851_ = ~new_n1176_ | ~new_n1528_;
  assign new_n1852_ = ~new_n1177_ | ~new_n1535_;
  assign new_n1853_ = ~new_n1178_ | ~new_n1263_;
  assign new_n1854_ = ~new_n1179_ | ~new_n1274_;
  assign new_n1855_ = ~new_n1180_ | ~new_n1532_;
  assign new_n1856_ = ~new_n1181_ | ~new_n1340_;
  assign new_n1857_ = ~new_n1182_ | ~new_n1276_;
  assign new_n1858_ = ~new_n1183_ | ~new_n1543_;
  assign new_n1859_ = ~new_n1188_ | ~new_n1538_;
  assign new_n1860_ = ~new_n1189_ | ~new_n1350_;
  assign new_n1861_ = ~new_n1192_ | ~new_n1552_;
  assign new_n1862_ = ~new_n1197_ | ~new_n1547_;
  assign new_n1863_ = ~new_n1200_ | ~new_n1568_;
  assign new_n1864_ = ~new_n1201_ | ~new_n1561_;
  assign new_n1865_ = ~new_n1206_ | ~new_n1556_;
  assign new_n1866_ = ~new_n1207_ | ~new_n1565_;
  assign new_n1867_ = ~new_n1210_ | ~new_n1562_;
  assign new_n1868_ = ~new_n1567_ | ~new_n1566_;
  assign new_n1869_ = ~new_n1213_ | ~new_n1555_;
  assign new_n1870_ = ~new_n1571_;
  assign new_n1871_ = ~new_n427_ | ~new_n1774_;
  assign new_n1872_ = ~new_n428_ | ~new_n1776_;
  assign new_n1873_ = ~new_n429_ | ~new_n1797_;
  assign new_n1874_ = ~new_n430_ | ~new_n1799_;
  assign new_n1875_ = ~new_n431_ | ~new_n1816_;
  assign new_n1876_ = ~new_n432_ | ~new_n1815_;
  assign new_n1877_ = ~new_n1578_;
  assign new_n1878_ = ~new_n1579_;
  assign new_n1879_ = ~new_n433_ | ~new_n1812_;
  assign new_n1880_ = ~new_n434_ | ~new_n1813_;
  assign new_n1881_ = ~new_n435_ | ~new_n1803_;
  assign new_n1882_ = ~new_n436_ | ~new_n1801_;
  assign new_n1883_ = ~new_n437_ | ~new_n1711_;
  assign new_n1884_ = ~new_n438_ | ~new_n1712_;
  assign new_n1885_ = ~new_n439_ | ~new_n1744_;
  assign new_n1886_ = ~new_n440_ | ~new_n1745_;
  assign new_n1887_ = ~new_n441_ | ~new_n1739_;
  assign new_n1888_ = ~new_n442_ | ~new_n1740_;
  assign new_n1889_ = ~new_n1592_;
  assign new_n1890_ = ~new_n443_ | ~new_n1721_;
  assign new_n1891_ = ~new_n444_ | ~new_n1722_;
  assign new_n1892_ = ~new_n445_ | ~new_n1734_;
  assign new_n1893_ = ~new_n446_ | ~new_n1735_;
  assign new_n1894_ = ~new_n447_ | ~new_n1705_;
  assign new_n1895_ = ~new_n448_ | ~new_n1706_;
  assign new_n1896_ = ~new_n449_ | ~new_n1701_;
  assign new_n1897_ = ~new_n450_ | ~new_n1702_;
  assign new_n1898_ = ~new_n1602_;
  assign new_n1899_ = ~new_n1603_;
  assign new_n1900_ = ~new_n451_ | ~new_n1698_;
  assign new_n1901_ = ~new_n452_ | ~new_n1697_;
  assign new_n1902_ = ~new_n453_ | ~new_n1732_;
  assign new_n1903_ = ~new_n454_ | ~new_n1731_;
  assign new_n1904_ = ~new_n455_ | ~new_n1827_;
  assign new_n1905_ = ~new_n456_ | ~new_n1826_;
  assign new_n1906_ = ~new_n457_ | ~new_n1824_;
  assign new_n1907_ = ~new_n458_ | ~new_n1823_;
  assign new_n1908_ = ~new_n459_ | ~new_n1819_;
  assign new_n1909_ = ~new_n460_ | ~new_n1818_;
  assign new_n1910_ = ~new_n1620_ | ~new_n1616_;
  assign new_n1911_ = ~new_n1849_ | ~new_n1617_;
  assign new_n1912_ = ~new_n1257_ | ~new_n1618_;
  assign new_n1913_ = ~new_n1258_ | ~new_n1619_;
  assign new_n1914_ = ~new_n1850_ | ~new_n1621_;
  assign new_n1915_ = ~new_n1261_ | ~new_n1622_;
  assign new_n1916_ = ~new_n1262_ | ~new_n1623_;
  assign new_n1917_ = ~new_n1853_ | ~new_n1624_;
  assign new_n1918_ = ~new_n1632_ | ~new_n1625_;
  assign new_n1919_ = ~new_n1265_ | ~new_n1626_;
  assign new_n1920_ = ~new_n1266_ | ~new_n1627_;
  assign new_n1921_ = ~new_n1269_ | ~new_n1630_;
  assign new_n1922_ = ~new_n1272_ | ~new_n1631_;
  assign new_n1923_ = ~new_n1854_ | ~new_n1633_;
  assign new_n1924_ = ~new_n1641_ | ~new_n1634_;
  assign new_n1925_ = ~new_n1857_ | ~new_n1635_;
  assign new_n1926_ = ~new_n1277_ | ~new_n1636_;
  assign new_n1927_ = ~new_n1278_ | ~new_n1637_;
  assign new_n1928_ = ~new_n1279_ | ~new_n1638_;
  assign new_n1929_ = ~new_n1280_ | ~new_n1639_;
  assign new_n1930_ = ~new_n1688_ | ~new_n1640_;
  assign new_n1931_ = ~new_n1649_ | ~new_n1642_;
  assign new_n1932_ = ~new_n1687_ | ~new_n1643_;
  assign new_n1933_ = ~new_n1285_ | ~new_n1644_;
  assign new_n1934_ = ~new_n1286_ | ~new_n1645_;
  assign new_n1935_ = ~new_n1287_ | ~new_n1646_;
  assign new_n1936_ = ~new_n1288_ | ~new_n1647_;
  assign new_n1937_ = ~new_n1684_ | ~new_n1648_;
  assign new_n1938_ = ~new_n1293_ | ~new_n1651_;
  assign new_n1939_ = ~new_n1654_ | ~new_n1294_;
  assign new_n1940_ = ~new_n1690_ | ~new_n1652_;
  assign new_n1941_ = ~new_n1297_ | ~new_n1653_;
  assign new_n1942_ = ~new_n1655_;
  assign new_n1943_ = ~new_n1656_;
  assign new_n1944_ = ~new_n1657_;
  assign new_n1945_ = ~new_n1659_ | ~new_n1663_;
  assign new_n1946_ = ~new_n1660_;
  assign new_n1947_ = ~new_n1661_ | ~new_n1662_;
  assign new_n1948_ = ~new_n1673_ | ~new_n1666_;
  assign new_n1949_ = ~new_n1847_ | ~new_n1667_;
  assign new_n1950_ = ~new_n1317_ | ~new_n1668_;
  assign new_n1951_ = ~new_n1318_ | ~new_n1669_;
  assign new_n1952_ = ~new_n1319_ | ~new_n1670_;
  assign new_n1953_ = ~new_n1320_ | ~new_n1671_;
  assign new_n1954_ = ~new_n1838_ | ~new_n1672_;
  assign new_n1955_ = ~new_n1323_ | ~new_n1674_;
  assign new_n1956_ = ~new_n1842_ | ~new_n1675_;
  assign new_n1957_ = ~new_n1676_ | ~new_n1725_;
  assign new_n1958_ = ~new_n1326_ | ~new_n1677_;
  assign new_n1959_ = ~new_n1329_ | ~new_n1679_;
  assign new_n1960_ = ~new_n1682_ | ~new_n1330_;
  assign new_n1961_ = ~new_n1844_ | ~new_n1680_;
  assign new_n1962_ = ~new_n1333_ | ~new_n1681_;
  assign new_n1963_ = ~new_n1683_ | ~new_n1334_;
  assign new_n1964_ = ~new_n1685_ | ~new_n1686_;
  assign new_n1965_ = ~new_n1689_ | ~new_n1856_;
  assign new_n1966_ = ~new_n1691_ | ~new_n1343_;
  assign new_n1967_ = ~new_n1692_ | ~new_n1693_;
  assign new_n1968_ = ~new_n1694_ | ~new_n1860_;
  assign new_n1969_ = ~new_n1356_ | ~new_n1704_;
  assign new_n1970_ = ~new_n1358_ | ~new_n1796_;
  assign new_n1971_ = ~new_n1361_ | ~new_n1700_;
  assign new_n1972_ = ~new_n1362_ | ~new_n1699_;
  assign new_n1973_ = ~new_n1366_ | ~new_n1794_;
  assign new_n1974_ = ~new_n1367_ | ~new_n1695_;
  assign new_n1975_ = ~new_n1370_ | ~new_n1733_;
  assign new_n1976_ = ~new_n1372_ | ~new_n1791_;
  assign new_n1977_ = ~new_n1373_ | ~new_n1737_;
  assign new_n1978_ = ~new_n1374_ | ~new_n1802_;
  assign new_n1979_ = ~new_n1378_ | ~new_n1748_;
  assign new_n1980_ = ~new_n1381_ | ~new_n1758_;
  assign new_n1981_ = ~new_n1087_ | ~new_n1718_;
  assign new_n1982_ = ~new_n1088_ | ~new_n1720_;
  assign new_n1983_ = ~new_n1388_ | ~new_n1723_;
  assign new_n1984_ = ~new_n1389_ | ~new_n1724_;
  assign new_n1985_ = ~new_n1840_ | ~new_n1726_;
  assign new_n1986_ = ~new_n1392_ | ~new_n1771_;
  assign new_n1987_ = ~new_n1395_ | ~new_n1828_;
  assign new_n1988_ = ~new_n1398_ | ~new_n1707_;
  assign new_n1989_ = ~new_n1401_ | ~new_n1790_;
  assign new_n1990_ = ~new_n1403_ | ~new_n1709_;
  assign new_n1991_ = ~new_n1404_ | ~new_n1743_;
  assign new_n1992_ = ~new_n1408_ | ~new_n1756_;
  assign new_n1993_ = ~new_n1409_ | ~new_n1747_;
  assign new_n1994_ = ~new_n1410_ | ~new_n1738_;
  assign new_n1995_ = ~new_n1413_ | ~new_n1787_;
  assign new_n1996_ = ~new_n1415_ | ~new_n1742_;
  assign new_n1997_ = ~new_n1416_ | ~new_n1713_;
  assign new_n1998_ = ~new_n1417_ | ~new_n1752_;
  assign new_n1999_ = ~new_n1419_ | ~new_n1749_;
  assign new_n2000_ = ~new_n1421_ | ~new_n1786_;
  assign new_n2001_ = ~new_n1422_ | ~new_n1741_;
  assign new_n2002_ = ~new_n1423_ | ~new_n1788_;
  assign new_n2003_ = ~new_n1424_ | ~new_n1716_;
  assign new_n2004_ = ~new_n1426_ | ~new_n1769_;
  assign new_n2005_ = ~new_n1429_ | ~new_n1770_;
  assign new_n2006_ = ~new_n1431_ | ~new_n1761_;
  assign new_n2007_ = ~new_n1432_ | ~new_n1766_;
  assign new_n2008_ = ~new_n1433_ | ~new_n1727_;
  assign new_n2009_ = ~new_n1773_ | ~new_n1772_;
  assign new_n2010_ = ~new_n1437_ | ~new_n1798_;
  assign new_n2011_ = ~new_n1800_ | ~new_n1777_;
  assign new_n2012_ = ~new_n1115_ | ~new_n1779_;
  assign new_n2013_ = ~new_n1443_ | ~new_n1783_;
  assign new_n2014_ = ~new_n1445_ | ~new_n1780_;
  assign new_n2015_ = ~new_n1447_ | ~new_n1755_;
  assign new_n2016_ = ~new_n1448_ | ~new_n1746_;
  assign new_n2017_ = ~new_n1449_ | ~new_n1757_;
  assign new_n2018_ = ~new_n1120_ | ~new_n1760_;
  assign new_n2019_ = ~new_n1451_ | ~new_n1792_;
  assign new_n2020_ = ~new_n1452_ | ~new_n1736_;
  assign new_n2021_ = ~new_n1453_ | ~new_n1708_;
  assign new_n2022_ = ~new_n1454_ | ~new_n1789_;
  assign new_n2023_ = ~new_n1455_ | ~new_n1795_;
  assign new_n2024_ = ~new_n1456_ | ~new_n1703_;
  assign new_n2025_ = ~new_n1457_ | ~new_n1793_;
  assign new_n2026_ = ~new_n1458_ | ~new_n1696_;
  assign new_n2027_ = ~new_n1460_ | ~new_n1775_;
  assign new_n2028_ = ~new_n1126_ | ~new_n1782_;
  assign new_n2029_ = ~new_n1128_ | ~new_n1751_;
  assign new_n2030_ = ~new_n1129_ | ~new_n1715_;
  assign new_n2031_ = ~new_n1469_ | ~new_n1710_;
  assign new_n2032_ = ~new_n1804_ | ~new_n1471_;
  assign new_n2033_ = ~new_n1132_ | ~new_n1806_;
  assign new_n2034_ = ~new_n1807_;
  assign new_n2035_ = ~new_n1657_ | ~new_n938_;
  assign new_n2036_ = ~new_n1477_ | ~new_n1808_;
  assign new_n2037_ = ~new_n1478_ | ~new_n1809_;
  assign new_n2038_ = ~new_n1656_ | ~new_n831_;
  assign new_n2039_ = ~new_n1141_ | ~new_n1754_;
  assign new_n2040_ = ~new_n1810_ | ~new_n1817_;
  assign new_n2041_ = ~new_n1482_ | ~new_n1814_;
  assign new_n2042_ = ~new_n1485_ | ~new_n1811_;
  assign new_n2043_ = ~new_n1145_ | ~new_n1785_;
  assign new_n2044_ = ~new_n1493_ | ~new_n1822_;
  assign new_n2045_ = ~new_n1148_ | ~new_n1768_;
  assign new_n2046_ = ~new_n1821_ | ~new_n1825_;
  assign new_n2047_ = ~new_n1497_ | ~new_n1820_;
  assign new_n2048_ = ~new_n1151_ | ~new_n1763_;
  assign new_n2049_ = ~new_n1505_ | ~new_n1730_;
  assign new_n2050_ = ~new_n1154_ | ~new_n1765_;
  assign new_n2051_ = ~new_n1155_ | ~new_n1729_;
  assign new_n2052_ = ~new_n1156_ | ~new_n1833_;
  assign new_n2053_ = new_n1831_;
  assign new_n2054_ = ~new_n1835_ | ~new_n1511_;
  assign new_n2055_ = ~new_n1832_;
  assign new_n2056_ = ~new_n1834_ | ~new_n1512_;
  assign new_n2057_ = ~new_n1834_;
  assign new_n2058_ = ~new_n1835_;
  assign new_n2059_ = ~new_n1836_ | ~new_n1843_;
  assign new_n2060_ = ~new_n1837_ | ~new_n1846_;
  assign new_n2061_ = ~new_n1841_ | ~new_n1839_;
  assign new_n2062_ = ~new_n1845_;
  assign new_n2063_ = ~new_n1851_ | ~new_n1848_;
  assign new_n2064_ = ~new_n1855_ | ~new_n1852_;
  assign new_n2065_ = ~new_n1859_ | ~new_n1858_;
  assign new_n2066_ = ~new_n1862_ | ~new_n1861_;
  assign new_n2067_ = ~new_n1863_ | ~new_n1869_;
  assign new_n2068_ = ~new_n1865_ | ~new_n1864_;
  assign new_n2069_ = ~new_n1867_ | ~new_n1866_;
  assign new_n2070_ = ~new_n1868_;
  assign new_n2071_ = ~new_n2034_ | ~new_n1870_;
  assign new_n2072_ = ~new_n1572_ | ~new_n1871_;
  assign new_n2073_ = ~new_n1573_ | ~new_n1872_;
  assign new_n2074_ = ~new_n1574_ | ~new_n1873_;
  assign new_n2075_ = ~new_n1575_ | ~new_n1874_;
  assign new_n2076_ = ~new_n1576_ | ~new_n1875_;
  assign new_n2077_ = ~new_n1577_ | ~new_n1876_;
  assign new_n2078_ = ~new_n1581_ | ~new_n1879_;
  assign new_n2079_ = ~new_n1582_ | ~new_n1880_;
  assign new_n2080_ = ~new_n1584_ | ~new_n1881_;
  assign new_n2081_ = ~new_n1585_ | ~new_n1882_;
  assign new_n2082_ = ~new_n1586_ | ~new_n1883_;
  assign new_n2083_ = ~new_n1587_ | ~new_n1884_;
  assign new_n2084_ = ~new_n1588_ | ~new_n1885_;
  assign new_n2085_ = ~new_n1589_ | ~new_n1886_;
  assign new_n2086_ = ~new_n1590_ | ~new_n1887_;
  assign new_n2087_ = ~new_n1591_ | ~new_n1888_;
  assign new_n2088_ = ~new_n1593_ | ~new_n1890_;
  assign new_n2089_ = ~new_n1595_ | ~new_n1891_;
  assign new_n2090_ = ~new_n1596_ | ~new_n1892_;
  assign new_n2091_ = ~new_n1597_ | ~new_n1893_;
  assign new_n2092_ = ~new_n1598_ | ~new_n1894_;
  assign new_n2093_ = ~new_n1599_ | ~new_n1895_;
  assign new_n2094_ = ~new_n1600_ | ~new_n1896_;
  assign new_n2095_ = ~new_n1601_ | ~new_n1897_;
  assign new_n2096_ = ~new_n1605_ | ~new_n1900_;
  assign new_n2097_ = ~new_n1606_ | ~new_n1901_;
  assign new_n2098_ = ~new_n1608_ | ~new_n1902_;
  assign new_n2099_ = ~new_n1609_ | ~new_n1903_;
  assign new_n2100_ = ~new_n1610_ | ~new_n1904_;
  assign new_n2101_ = ~new_n1611_ | ~new_n1905_;
  assign new_n2102_ = ~new_n1612_ | ~new_n1906_;
  assign new_n2103_ = ~new_n1613_ | ~new_n1907_;
  assign new_n2104_ = ~new_n1614_ | ~new_n1908_;
  assign new_n2105_ = ~new_n1615_ | ~new_n1909_;
  assign new_n2106_ = ~new_n1910_;
  assign new_n2107_ = new_n1911_ & new_n1914_ & new_n1923_ & new_n1917_;
  assign new_n2108_ = new_n1912_ & new_n1916_ & new_n1922_ & new_n1919_;
  assign new_n2109_ = new_n1912_;
  assign new_n2110_ = new_n1912_;
  assign new_n2111_ = new_n1913_;
  assign new_n2112_ = new_n1913_;
  assign new_n2113_ = new_n1913_ & new_n1920_ & new_n1915_ & new_n1921_;
  assign new_n2114_ = new_n1911_ & new_n981_;
  assign new_n2115_ = new_n1913_ & new_n984_;
  assign new_n2116_ = new_n1915_;
  assign new_n2117_ = new_n1915_;
  assign new_n2118_ = new_n1915_ & new_n1921_ & new_n1920_;
  assign new_n2119_ = new_n1912_ & new_n985_;
  assign new_n2120_ = new_n1916_;
  assign new_n2121_ = new_n1916_ & new_n1922_ & new_n1919_;
  assign new_n2122_ = new_n1916_;
  assign new_n2123_ = new_n1916_ & new_n986_;
  assign new_n2124_ = new_n986_ & new_n1916_ & new_n1912_;
  assign new_n2125_ = new_n1916_ & new_n986_;
  assign new_n2126_ = new_n987_ & new_n1915_ & new_n1913_;
  assign new_n2127_ = new_n1915_ & new_n987_;
  assign new_n2128_ = new_n1915_ & new_n987_;
  assign new_n2129_ = new_n988_ & new_n1914_ & new_n1911_;
  assign new_n2130_ = ~new_n1918_;
  assign new_n2131_ = new_n1922_ & new_n1919_;
  assign new_n2132_ = new_n1919_;
  assign new_n2133_ = new_n1919_;
  assign new_n2134_ = new_n1920_;
  assign new_n2135_ = new_n1920_;
  assign new_n2136_ = new_n1921_ & new_n1920_;
  assign new_n2137_ = new_n1916_ & new_n1919_ & new_n991_;
  assign new_n2138_ = new_n1916_ & new_n991_ & new_n1919_ & new_n1912_;
  assign new_n2139_ = new_n1916_ & new_n1919_ & new_n991_;
  assign new_n2140_ = new_n1919_ & new_n991_;
  assign new_n2141_ = new_n1915_ & new_n992_ & new_n1920_ & new_n1913_;
  assign new_n2142_ = new_n1915_ & new_n992_ & new_n1920_;
  assign new_n2143_ = new_n1915_ & new_n1920_ & new_n992_;
  assign new_n2144_ = new_n1920_ & new_n992_;
  assign new_n2145_ = new_n1920_ & new_n992_;
  assign new_n2146_ = ~new_n1921_;
  assign new_n2147_ = new_n1922_;
  assign new_n2148_ = new_n1922_;
  assign new_n2149_ = new_n1914_ & new_n995_ & new_n1917_ & new_n1911_;
  assign new_n2150_ = new_n1924_;
  assign new_n2151_ = new_n1924_;
  assign new_n2152_ = new_n1925_ & new_n1930_ & new_n1932_ & new_n1940_ & new_n1937_;
  assign new_n2153_ = new_n1926_;
  assign new_n2154_ = new_n1926_;
  assign new_n2155_ = new_n1926_ & new_n1929_ & new_n1933_ & new_n1938_ & new_n1936_;
  assign new_n2156_ = new_n1935_ & new_n1927_ & new_n1934_ & new_n1928_ & new_n1941_;
  assign new_n2157_ = new_n1927_;
  assign new_n2158_ = new_n1926_ & new_n1003_;
  assign new_n2159_ = new_n1927_ & new_n1004_;
  assign new_n2160_ = new_n1928_;
  assign new_n2161_ = new_n1929_;
  assign new_n2162_ = new_n1936_ & new_n1929_ & new_n1938_ & new_n1933_;
  assign new_n2163_ = new_n1929_;
  assign new_n2164_ = new_n1925_ & new_n1005_;
  assign new_n2165_ = new_n1929_ & new_n1008_;
  assign new_n2166_ = new_n1929_ & new_n1008_;
  assign new_n2167_ = new_n1008_ & new_n1929_ & new_n1926_;
  assign new_n2168_ = new_n1928_ & new_n1009_;
  assign new_n2169_ = new_n1009_ & new_n1928_ & new_n1927_;
  assign new_n2170_ = new_n1010_ & new_n1930_ & new_n1925_;
  assign new_n2171_ = ~new_n1931_;
  assign new_n2172_ = new_n1933_;
  assign new_n2173_ = new_n1933_;
  assign new_n2174_ = new_n1936_ & new_n1938_ & new_n1933_;
  assign new_n2175_ = new_n1934_;
  assign new_n2176_ = new_n1929_ & new_n1933_ & new_n1013_;
  assign new_n2177_ = new_n1929_ & new_n1933_ & new_n1013_;
  assign new_n2178_ = new_n1929_ & new_n1013_ & new_n1933_ & new_n1926_;
  assign new_n2179_ = new_n1933_ & new_n1013_;
  assign new_n2180_ = new_n1933_ & new_n1013_;
  assign new_n2181_ = new_n1928_ & new_n1934_ & new_n1014_;
  assign new_n2182_ = new_n1928_ & new_n1014_ & new_n1934_ & new_n1927_;
  assign new_n2183_ = new_n1014_ & new_n1934_;
  assign new_n2184_ = new_n1935_;
  assign new_n2185_ = new_n1936_;
  assign new_n2186_ = new_n1936_;
  assign new_n2187_ = new_n1938_ & new_n1936_;
  assign new_n2188_ = new_n1930_ & new_n1015_ & new_n1932_ & new_n1925_;
  assign new_n2189_ = new_n1929_ & new_n1018_ & new_n1936_ & new_n1933_;
  assign new_n2190_ = new_n1929_ & new_n1018_ & new_n1926_ & new_n1936_ & new_n1933_;
  assign new_n2191_ = new_n1929_ & new_n1018_ & new_n1936_ & new_n1933_;
  assign new_n2192_ = new_n1018_ & new_n1936_ & new_n1933_;
  assign new_n2193_ = new_n1936_ & new_n1018_;
  assign new_n2194_ = new_n1018_ & new_n1936_ & new_n1933_;
  assign new_n2195_ = new_n1928_ & new_n1019_ & new_n1935_ & new_n1934_;
  assign new_n2196_ = new_n1928_ & new_n1019_ & new_n1927_ & new_n1935_ & new_n1934_;
  assign new_n2197_ = new_n1935_ & new_n1019_;
  assign new_n2198_ = new_n1019_ & new_n1935_ & new_n1934_;
  assign new_n2199_ = new_n1938_;
  assign new_n2200_ = new_n1938_;
  assign new_n2201_ = new_n1930_ & new_n1021_ & new_n1925_ & new_n1937_ & new_n1932_;
  assign new_n2202_ = ~new_n1939_;
  assign new_n2203_ = new_n1941_;
  assign new_n2204_ = new_n1948_;
  assign new_n2205_ = new_n1948_;
  assign new_n2206_ = new_n1949_ & new_n1954_ & new_n1985_ & new_n1961_ & new_n1956_;
  assign new_n2207_ = new_n1950_;
  assign new_n2208_ = new_n1950_;
  assign new_n2209_ = new_n1950_ & new_n1953_ & new_n1983_ & new_n1959_ & new_n1958_;
  assign new_n2210_ = new_n1955_ & new_n1951_ & new_n1984_ & new_n1952_ & new_n1962_;
  assign new_n2211_ = new_n1951_;
  assign new_n2212_ = new_n1950_ & new_n1038_;
  assign new_n2213_ = new_n1951_ & new_n1039_;
  assign new_n2214_ = new_n1952_;
  assign new_n2215_ = new_n1953_;
  assign new_n2216_ = new_n1958_ & new_n1953_ & new_n1959_ & new_n1983_;
  assign new_n2217_ = new_n1953_;
  assign new_n2218_ = new_n1949_ & new_n1040_;
  assign new_n2219_ = new_n1953_ & new_n1983_ & new_n1043_;
  assign new_n2220_ = new_n1953_ & new_n1983_ & new_n1043_;
  assign new_n2221_ = new_n1953_ & new_n1043_ & new_n1983_ & new_n1950_;
  assign new_n2222_ = new_n1983_ & new_n1043_;
  assign new_n2223_ = new_n1983_ & new_n1043_;
  assign new_n2224_ = new_n1952_ & new_n1984_ & new_n1044_;
  assign new_n2225_ = new_n1952_ & new_n1044_ & new_n1984_ & new_n1951_;
  assign new_n2226_ = new_n1044_ & new_n1984_;
  assign new_n2227_ = new_n1955_;
  assign new_n2228_ = new_n1954_ & new_n1045_ & new_n1985_ & new_n1949_;
  assign new_n2229_ = ~new_n1957_;
  assign new_n2230_ = new_n1958_;
  assign new_n2231_ = new_n1958_ & new_n1959_ & new_n1983_;
  assign new_n2232_ = new_n1958_;
  assign new_n2233_ = new_n1959_ & new_n1958_;
  assign new_n2234_ = new_n1953_ & new_n1048_ & new_n1958_ & new_n1983_;
  assign new_n2235_ = new_n1953_ & new_n1048_ & new_n1950_ & new_n1958_ & new_n1983_;
  assign new_n2236_ = new_n1953_ & new_n1048_ & new_n1958_ & new_n1983_;
  assign new_n2237_ = new_n1048_ & new_n1958_ & new_n1983_;
  assign new_n2238_ = new_n1958_ & new_n1048_;
  assign new_n2239_ = new_n1048_ & new_n1958_ & new_n1983_;
  assign new_n2240_ = new_n1952_ & new_n1049_ & new_n1955_ & new_n1984_;
  assign new_n2241_ = new_n1952_ & new_n1049_ & new_n1951_ & new_n1955_ & new_n1984_;
  assign new_n2242_ = new_n1955_ & new_n1049_;
  assign new_n2243_ = new_n1049_ & new_n1955_ & new_n1984_;
  assign new_n2244_ = new_n1959_;
  assign new_n2245_ = new_n1959_;
  assign new_n2246_ = new_n1954_ & new_n1051_ & new_n1949_ & new_n1956_ & new_n1985_;
  assign new_n2247_ = ~new_n1960_;
  assign new_n2248_ = new_n1962_;
  assign new_n2249_ = ~new_n1963_;
  assign new_n2250_ = ~new_n1964_;
  assign new_n2251_ = new_n1965_;
  assign new_n2252_ = new_n1965_;
  assign new_n2253_ = ~new_n1966_;
  assign new_n2254_ = ~new_n1967_;
  assign new_n2255_ = new_n1968_;
  assign new_n2256_ = new_n1968_;
  assign new_n2257_ = ~new_n1969_ | ~new_n1974_;
  assign new_n2258_ = ~new_n1970_ | ~new_n2026_;
  assign new_n2259_ = ~new_n1971_ | ~new_n1972_;
  assign new_n2260_ = ~new_n1973_ | ~new_n2024_;
  assign new_n2261_ = ~new_n1975_ | ~new_n1988_;
  assign new_n2262_ = ~new_n1976_ | ~new_n2021_;
  assign new_n2263_ = ~new_n1977_ | ~new_n1990_;
  assign new_n2264_ = ~new_n1978_ | ~new_n2031_;
  assign new_n2265_ = ~new_n1979_ | ~new_n1997_;
  assign new_n2266_ = ~new_n1714_ | ~new_n2030_;
  assign new_n2267_ = ~new_n1980_ | ~new_n2003_;
  assign new_n2268_ = ~new_n1981_ | ~new_n1717_;
  assign new_n2269_ = ~new_n1982_ | ~new_n1719_;
  assign new_n2270_ = new_n1953_ & new_n1089_;
  assign new_n2271_ = new_n1953_ & new_n1089_;
  assign new_n2272_ = new_n1089_ & new_n1953_ & new_n1950_;
  assign new_n2273_ = new_n1952_ & new_n1090_;
  assign new_n2274_ = new_n1090_ & new_n1952_ & new_n1951_;
  assign new_n2275_ = new_n1983_;
  assign new_n2276_ = new_n1983_;
  assign new_n2277_ = new_n1984_;
  assign new_n2278_ = new_n1091_ & new_n1954_ & new_n1949_;
  assign new_n2279_ = ~new_n1986_ | ~new_n2008_;
  assign new_n2280_ = ~new_n2051_ | ~new_n1728_;
  assign new_n2281_ = ~new_n2049_ | ~new_n1987_;
  assign new_n2282_ = ~new_n1989_ | ~new_n2020_;
  assign new_n2283_ = ~new_n1991_ | ~new_n1994_;
  assign new_n2284_ = ~new_n1992_ | ~new_n2001_;
  assign new_n2285_ = ~new_n1993_ | ~new_n1996_;
  assign new_n2286_ = ~new_n1995_ | ~new_n2016_;
  assign new_n2287_ = ~new_n1998_ | ~new_n1999_;
  assign new_n2288_ = ~new_n2029_ | ~new_n1750_;
  assign new_n2289_ = ~new_n2039_ | ~new_n1753_;
  assign new_n2290_ = ~new_n2000_ | ~new_n2015_;
  assign new_n2291_ = ~new_n2002_ | ~new_n2017_;
  assign new_n2292_ = ~new_n2018_ | ~new_n1759_;
  assign new_n2293_ = ~new_n2006_ | ~new_n2004_;
  assign new_n2294_ = ~new_n2048_ | ~new_n1762_;
  assign new_n2295_ = ~new_n2050_ | ~new_n1764_;
  assign new_n2296_ = ~new_n2005_ | ~new_n2007_;
  assign new_n2297_ = ~new_n2045_ | ~new_n1767_;
  assign new_n2298_ = ~new_n2009_;
  assign new_n2299_ = ~new_n2027_ | ~new_n2010_;
  assign new_n2300_ = ~new_n2011_;
  assign new_n2301_ = ~new_n2012_ | ~new_n1778_;
  assign new_n2302_ = ~new_n2014_ | ~new_n2013_;
  assign new_n2303_ = ~new_n2028_ | ~new_n1781_;
  assign new_n2304_ = ~new_n2043_ | ~new_n1784_;
  assign new_n2305_ = ~new_n2022_ | ~new_n2019_;
  assign new_n2306_ = ~new_n2025_ | ~new_n2023_;
  assign new_n2307_ = ~new_n2032_;
  assign new_n2308_ = ~new_n2033_ | ~new_n1805_;
  assign new_n2309_ = ~new_n827_ | ~new_n1944_;
  assign new_n2310_ = ~new_n2037_;
  assign new_n2311_ = ~new_n673_ | ~new_n1943_;
  assign new_n2312_ = ~new_n2040_;
  assign new_n2313_ = ~new_n2041_ | ~new_n2042_;
  assign new_n2314_ = ~new_n2044_ | ~new_n2047_;
  assign new_n2315_ = ~new_n2046_;
  assign new_n2316_ = ~new_n1829_ | ~new_n2052_;
  assign new_n2317_ = ~new_n2053_;
  assign new_n2318_ = ~new_n1157_ | ~new_n2058_;
  assign new_n2319_ = ~new_n1158_ | ~new_n2057_;
  assign new_n2320_ = ~new_n2059_;
  assign new_n2321_ = new_n2060_;
  assign new_n2322_ = new_n2060_;
  assign new_n2323_ = ~new_n2061_;
  assign new_n2324_ = ~new_n2063_;
  assign new_n2325_ = ~new_n2064_;
  assign new_n2326_ = ~new_n2065_;
  assign new_n2327_ = ~new_n2066_;
  assign new_n2328_ = new_n2067_;
  assign new_n2329_ = new_n2067_;
  assign new_n2330_ = ~new_n2068_;
  assign new_n2331_ = ~new_n2069_;
  assign new_n2332_ = new_n1571_ & new_n2206_;
  assign new_n2333_ = new_n2072_ & new_n2075_ & new_n2078_ & new_n2077_;
  assign new_n2334_ = new_n2072_;
  assign new_n2335_ = new_n2072_;
  assign new_n2336_ = new_n2073_;
  assign new_n2337_ = new_n2073_;
  assign new_n2338_ = new_n2073_ & new_n2076_ & new_n2074_ & new_n2079_;
  assign new_n2339_ = new_n2073_ & new_n1218_;
  assign new_n2340_ = new_n2072_ & new_n1219_;
  assign new_n2341_ = new_n2074_;
  assign new_n2342_ = new_n2074_;
  assign new_n2343_ = new_n2074_ & new_n2079_ & new_n2076_;
  assign new_n2344_ = new_n2075_;
  assign new_n2345_ = new_n2075_ & new_n2078_ & new_n2077_;
  assign new_n2346_ = new_n2075_;
  assign new_n2347_ = new_n1220_ & new_n2074_ & new_n2073_;
  assign new_n2348_ = new_n2074_ & new_n1220_;
  assign new_n2349_ = new_n2074_ & new_n1220_;
  assign new_n2350_ = new_n2075_ & new_n1221_;
  assign new_n2351_ = new_n1221_ & new_n2075_ & new_n2072_;
  assign new_n2352_ = new_n2075_ & new_n1221_;
  assign new_n2353_ = new_n2076_;
  assign new_n2354_ = new_n2076_;
  assign new_n2355_ = new_n2079_ & new_n2076_;
  assign new_n2356_ = new_n2078_ & new_n2077_;
  assign new_n2357_ = new_n2077_;
  assign new_n2358_ = new_n2077_;
  assign new_n2359_ = new_n2074_ & new_n1222_ & new_n2076_ & new_n2073_;
  assign new_n2360_ = new_n2074_ & new_n1222_ & new_n2076_;
  assign new_n2361_ = new_n2074_ & new_n2076_ & new_n1222_;
  assign new_n2362_ = new_n2076_ & new_n1222_;
  assign new_n2363_ = new_n2076_ & new_n1222_;
  assign new_n2364_ = new_n2075_ & new_n2077_ & new_n1223_;
  assign new_n2365_ = new_n2075_ & new_n1223_ & new_n2077_ & new_n2072_;
  assign new_n2366_ = new_n2075_ & new_n2077_ & new_n1223_;
  assign new_n2367_ = new_n2077_ & new_n1223_;
  assign new_n2368_ = new_n2078_;
  assign new_n2369_ = new_n2078_;
  assign new_n2370_ = ~new_n2079_;
  assign new_n2371_ = new_n2080_;
  assign new_n2372_ = new_n2080_;
  assign new_n2373_ = new_n2080_ & new_n2083_ & new_n2084_ & new_n2089_ & new_n2086_;
  assign new_n2374_ = new_n2087_ & new_n2081_ & new_n2085_ & new_n2082_ & new_n2088_;
  assign new_n2375_ = new_n2081_;
  assign new_n2376_ = new_n2081_ & new_n1228_;
  assign new_n2377_ = new_n2080_ & new_n1229_;
  assign new_n2378_ = new_n2082_;
  assign new_n2379_ = new_n2083_;
  assign new_n2380_ = new_n2086_ & new_n2083_ & new_n2089_ & new_n2084_;
  assign new_n2381_ = new_n2083_;
  assign new_n2382_ = new_n2082_ & new_n1230_;
  assign new_n2383_ = new_n1230_ & new_n2082_ & new_n2081_;
  assign new_n2384_ = new_n2083_ & new_n1231_;
  assign new_n2385_ = new_n2083_ & new_n1231_;
  assign new_n2386_ = new_n1231_ & new_n2083_ & new_n2080_;
  assign new_n2387_ = new_n2084_;
  assign new_n2388_ = new_n2084_;
  assign new_n2389_ = new_n2086_ & new_n2089_ & new_n2084_;
  assign new_n2390_ = new_n2085_;
  assign new_n2391_ = new_n2082_ & new_n2085_ & new_n1232_;
  assign new_n2392_ = new_n2082_ & new_n1232_ & new_n2085_ & new_n2081_;
  assign new_n2393_ = new_n1232_ & new_n2085_;
  assign new_n2394_ = new_n2083_ & new_n2084_ & new_n1233_;
  assign new_n2395_ = new_n2083_ & new_n2084_ & new_n1233_;
  assign new_n2396_ = new_n2083_ & new_n1233_ & new_n2084_ & new_n2080_;
  assign new_n2397_ = new_n2084_ & new_n1233_;
  assign new_n2398_ = new_n2084_ & new_n1233_;
  assign new_n2399_ = new_n2086_;
  assign new_n2400_ = new_n2086_;
  assign new_n2401_ = new_n2089_ & new_n2086_;
  assign new_n2402_ = new_n2087_;
  assign new_n2403_ = new_n2082_ & new_n1234_ & new_n2087_ & new_n2085_;
  assign new_n2404_ = new_n2082_ & new_n1234_ & new_n2081_ & new_n2087_ & new_n2085_;
  assign new_n2405_ = new_n2087_ & new_n1234_;
  assign new_n2406_ = new_n1234_ & new_n2087_ & new_n2085_;
  assign new_n2407_ = new_n2083_ & new_n1235_ & new_n2086_ & new_n2084_;
  assign new_n2408_ = new_n2083_ & new_n1235_ & new_n2080_ & new_n2086_ & new_n2084_;
  assign new_n2409_ = new_n2083_ & new_n1235_ & new_n2086_ & new_n2084_;
  assign new_n2410_ = new_n1235_ & new_n2086_ & new_n2084_;
  assign new_n2411_ = new_n2086_ & new_n1235_;
  assign new_n2412_ = new_n1235_ & new_n2086_ & new_n2084_;
  assign new_n2413_ = new_n2088_;
  assign new_n2414_ = new_n2089_;
  assign new_n2415_ = new_n2089_;
  assign new_n2416_ = new_n2090_ & new_n2093_ & new_n2096_ & new_n2094_;
  assign new_n2417_ = new_n2090_;
  assign new_n2418_ = new_n2090_;
  assign new_n2419_ = new_n2091_;
  assign new_n2420_ = new_n2091_;
  assign new_n2421_ = new_n2091_ & new_n2095_ & new_n2092_ & new_n2097_;
  assign new_n2422_ = new_n2091_ & new_n1239_;
  assign new_n2423_ = new_n2090_ & new_n1240_;
  assign new_n2424_ = new_n2092_;
  assign new_n2425_ = new_n2092_;
  assign new_n2426_ = new_n2092_ & new_n2097_ & new_n2095_;
  assign new_n2427_ = new_n2093_;
  assign new_n2428_ = new_n2093_ & new_n2096_ & new_n2094_;
  assign new_n2429_ = new_n2093_;
  assign new_n2430_ = new_n1241_ & new_n2092_ & new_n2091_;
  assign new_n2431_ = new_n2092_ & new_n1241_;
  assign new_n2432_ = new_n2092_ & new_n1241_;
  assign new_n2433_ = new_n2093_ & new_n1242_;
  assign new_n2434_ = new_n1242_ & new_n2093_ & new_n2090_;
  assign new_n2435_ = new_n2093_ & new_n1242_;
  assign new_n2436_ = new_n2096_ & new_n2094_;
  assign new_n2437_ = new_n2094_;
  assign new_n2438_ = new_n2094_;
  assign new_n2439_ = new_n2095_;
  assign new_n2440_ = new_n2095_;
  assign new_n2441_ = new_n2097_ & new_n2095_;
  assign new_n2442_ = new_n2092_ & new_n1243_ & new_n2095_ & new_n2091_;
  assign new_n2443_ = new_n2092_ & new_n1243_ & new_n2095_;
  assign new_n2444_ = new_n2092_ & new_n2095_ & new_n1243_;
  assign new_n2445_ = new_n2095_ & new_n1243_;
  assign new_n2446_ = new_n2095_ & new_n1243_;
  assign new_n2447_ = new_n2093_ & new_n2094_ & new_n1244_;
  assign new_n2448_ = new_n2093_ & new_n1244_ & new_n2094_ & new_n2090_;
  assign new_n2449_ = new_n2093_ & new_n2094_ & new_n1244_;
  assign new_n2450_ = new_n2094_ & new_n1244_;
  assign new_n2451_ = new_n2096_;
  assign new_n2452_ = new_n2096_;
  assign new_n2453_ = ~new_n2097_;
  assign new_n2454_ = new_n2098_;
  assign new_n2455_ = new_n2099_;
  assign new_n2456_ = new_n2099_;
  assign new_n2457_ = new_n2098_ & new_n1249_;
  assign new_n2458_ = new_n2099_ & new_n1250_;
  assign new_n2459_ = new_n2100_;
  assign new_n2460_ = new_n2100_;
  assign new_n2461_ = new_n2101_;
  assign new_n2462_ = new_n2101_ & new_n1251_;
  assign new_n2463_ = new_n1251_ & new_n2101_ & new_n2098_;
  assign new_n2464_ = new_n2100_ & new_n1252_;
  assign new_n2465_ = new_n2100_ & new_n1252_;
  assign new_n2466_ = new_n1252_ & new_n2100_ & new_n2099_;
  assign new_n2467_ = new_n2102_;
  assign new_n2468_ = new_n2103_;
  assign new_n2469_ = new_n2103_;
  assign new_n2470_ = new_n2101_ & new_n2102_ & new_n1253_;
  assign new_n2471_ = new_n2101_ & new_n1253_ & new_n2102_ & new_n2098_;
  assign new_n2472_ = new_n1253_ & new_n2102_;
  assign new_n2473_ = new_n2100_ & new_n2103_ & new_n1254_;
  assign new_n2474_ = new_n2100_ & new_n2103_ & new_n1254_;
  assign new_n2475_ = new_n2100_ & new_n1254_ & new_n2103_ & new_n2099_;
  assign new_n2476_ = new_n2103_ & new_n1254_;
  assign new_n2477_ = new_n2103_ & new_n1254_;
  assign new_n2478_ = new_n2104_;
  assign new_n2479_ = new_n2104_;
  assign new_n2480_ = new_n2105_;
  assign new_n2481_ = new_n2149_ | new_n2129_ | new_n976_ | new_n2114_;
  assign new_n2482_ = ~new_n1910_ | ~new_n2130_;
  assign new_n2483_ = new_n2107_ & new_n2152_;
  assign new_n2484_ = new_n2108_ & new_n2155_;
  assign new_n2485_ = ~new_n2109_;
  assign new_n2486_ = ~new_n2110_;
  assign new_n2487_ = new_n2138_ | new_n2124_ | new_n979_ | new_n2119_;
  assign new_n2488_ = new_n2141_ | new_n2126_ | new_n980_ | new_n2115_;
  assign new_n2489_ = ~new_n2111_;
  assign new_n2490_ = ~new_n2112_;
  assign new_n2491_ = new_n2113_ & new_n2156_;
  assign new_n2492_ = ~new_n2142_ & ~new_n984_ & ~new_n2128_;
  assign new_n2493_ = new_n2118_ | new_n2143_ | new_n984_ | new_n2127_;
  assign new_n2494_ = ~new_n2116_;
  assign new_n2495_ = ~new_n2117_;
  assign new_n2496_ = ~new_n2139_ & ~new_n985_ & ~new_n2123_;
  assign new_n2497_ = new_n2121_ | new_n2137_ | new_n985_ | new_n2125_;
  assign new_n2498_ = ~new_n2120_;
  assign new_n2499_ = ~new_n2122_;
  assign new_n2500_ = new_n986_ | new_n2140_;
  assign new_n2501_ = ~new_n987_ & ~new_n2145_;
  assign new_n2502_ = new_n2136_ | new_n987_ | new_n2144_;
  assign new_n2503_ = ~new_n1918_ | ~new_n2106_;
  assign new_n2504_ = ~new_n2132_;
  assign new_n2505_ = ~new_n2133_;
  assign new_n2506_ = ~new_n2134_;
  assign new_n2507_ = ~new_n2135_;
  assign new_n2508_ = ~new_n2134_ | ~new_n1629_;
  assign new_n2509_ = ~new_n2135_ | ~new_n1270_;
  assign new_n2510_ = ~new_n2147_;
  assign new_n2511_ = ~new_n2148_;
  assign new_n2512_ = new_n2201_ | new_n2188_ | new_n2170_ | new_n998_ | new_n2164_;
  assign new_n2513_ = new_n2150_ & new_n2171_ & new_n2202_;
  assign new_n2514_ = ~new_n2150_;
  assign new_n2515_ = ~new_n2151_;
  assign new_n2516_ = new_n2190_ | new_n2178_ | new_n2167_ | new_n1001_ | new_n2158_;
  assign new_n2517_ = ~new_n2153_;
  assign new_n2518_ = ~new_n2154_;
  assign new_n2519_ = ~new_n2155_;
  assign new_n2520_ = new_n2196_ | new_n2182_ | new_n2169_ | new_n1002_ | new_n2159_;
  assign new_n2521_ = ~new_n2157_;
  assign new_n2522_ = ~new_n2191_ & ~new_n2176_ & ~new_n1003_ & ~new_n2165_;
  assign new_n2523_ = new_n2162_ | new_n2189_ | new_n2177_ | new_n1003_ | new_n2166_;
  assign new_n2524_ = ~new_n2160_;
  assign new_n2525_ = ~new_n2161_;
  assign new_n2526_ = ~new_n2163_;
  assign new_n2527_ = ~new_n2194_ & ~new_n1008_ & ~new_n2179_;
  assign new_n2528_ = new_n2174_ | new_n2192_ | new_n1008_ | new_n2180_;
  assign new_n2529_ = new_n2151_ & new_n1931_ & new_n1939_;
  assign new_n2530_ = ~new_n2172_;
  assign new_n2531_ = ~new_n2173_;
  assign new_n2532_ = ~new_n2175_;
  assign new_n2533_ = new_n1013_ | new_n2193_;
  assign new_n2534_ = ~new_n2184_;
  assign new_n2535_ = ~new_n2185_;
  assign new_n2536_ = ~new_n2186_;
  assign new_n2537_ = ~new_n2199_;
  assign new_n2538_ = ~new_n2200_;
  assign new_n2539_ = ~new_n2203_;
  assign new_n2540_ = new_n1305_ & new_n2210_;
  assign new_n2541_ = new_n1308_ & new_n2209_;
  assign new_n2542_ = new_n2235_ | new_n2221_ | new_n2272_ | new_n1033_ | new_n2212_;
  assign new_n2543_ = new_n2241_ | new_n2225_ | new_n2274_ | new_n1034_ | new_n2213_;
  assign new_n2544_ = new_n2246_ | new_n2228_ | new_n2278_ | new_n1035_ | new_n2218_;
  assign new_n2545_ = new_n2204_ & new_n2229_ & new_n2247_;
  assign new_n2546_ = ~new_n2204_;
  assign new_n2547_ = ~new_n2205_;
  assign new_n2548_ = ~new_n2207_;
  assign new_n2549_ = ~new_n2208_;
  assign new_n2550_ = ~new_n2209_;
  assign new_n2551_ = ~new_n2211_;
  assign new_n2552_ = ~new_n2236_ & ~new_n2219_ & ~new_n1038_ & ~new_n2270_;
  assign new_n2553_ = new_n2216_ | new_n2234_ | new_n2220_ | new_n1038_ | new_n2271_;
  assign new_n2554_ = ~new_n2214_;
  assign new_n2555_ = ~new_n2215_;
  assign new_n2556_ = ~new_n2217_;
  assign new_n2557_ = new_n1043_ | new_n2238_;
  assign new_n2558_ = ~new_n2227_;
  assign new_n2559_ = new_n2205_ & new_n1957_ & new_n1960_;
  assign new_n2560_ = ~new_n2230_;
  assign new_n2561_ = ~new_n2232_;
  assign new_n2562_ = ~new_n2244_;
  assign new_n2563_ = ~new_n2245_;
  assign new_n2564_ = ~new_n2248_;
  assign new_n2565_ = new_n2251_ & new_n1964_ & new_n1963_;
  assign new_n2566_ = new_n2252_ & new_n2250_ & new_n2249_;
  assign new_n2567_ = ~new_n2251_;
  assign new_n2568_ = ~new_n2252_;
  assign new_n2569_ = new_n2255_ & new_n1967_ & new_n1966_;
  assign new_n2570_ = new_n2256_ & new_n2254_ & new_n2253_;
  assign new_n2571_ = ~new_n2255_;
  assign new_n2572_ = ~new_n2256_;
  assign new_n2573_ = ~new_n2257_;
  assign new_n2574_ = new_n2262_ & new_n1357_ & new_n2260_ & new_n2282_;
  assign new_n2575_ = new_n2282_ & new_n2262_ & new_n2258_ & new_n2260_;
  assign new_n2576_ = ~new_n2259_;
  assign new_n2577_ = new_n1365_ & new_n2262_ & new_n2282_;
  assign new_n2578_ = ~new_n2261_;
  assign new_n2579_ = new_n2282_ & new_n1371_;
  assign new_n2580_ = ~new_n2263_;
  assign new_n2581_ = new_n2264_;
  assign new_n2582_ = new_n2264_;
  assign new_n2583_ = new_n2288_ & new_n1377_;
  assign new_n2584_ = new_n2288_ & new_n2265_ & new_n2286_ & new_n2267_ & new_n2284_;
  assign new_n2585_ = new_n2266_;
  assign new_n2586_ = new_n2266_;
  assign new_n2587_ = new_n2265_ & new_n1380_ & new_n2288_ & new_n2284_ & new_n2286_;
  assign new_n2588_ = ~new_n2268_;
  assign new_n2589_ = ~new_n2269_;
  assign new_n2590_ = ~new_n2239_ & ~new_n1089_ & ~new_n2222_;
  assign new_n2591_ = new_n2231_ | new_n2237_ | new_n1089_ | new_n2223_;
  assign new_n2592_ = ~new_n2275_;
  assign new_n2593_ = ~new_n2276_;
  assign new_n2594_ = ~new_n2277_;
  assign new_n2595_ = new_n2279_ & new_n2295_ & new_n2294_ & new_n2316_ & new_n2297_;
  assign new_n2596_ = new_n2280_;
  assign new_n2597_ = new_n2280_;
  assign new_n2598_ = new_n2281_;
  assign new_n2599_ = new_n2281_;
  assign new_n2600_ = ~new_n2283_;
  assign new_n2601_ = new_n2265_ & new_n1407_ & new_n2286_ & new_n2288_;
  assign new_n2602_ = ~new_n2285_;
  assign new_n2603_ = new_n1414_ & new_n2265_ & new_n2288_;
  assign new_n2604_ = new_n2287_;
  assign new_n2605_ = new_n2287_;
  assign new_n2606_ = new_n2301_ & new_n2303_ & new_n2289_ & new_n2304_;
  assign new_n2607_ = ~new_n2290_;
  assign new_n2608_ = ~new_n2291_;
  assign new_n2609_ = ~new_n2292_;
  assign new_n2610_ = ~new_n2293_;
  assign new_n2611_ = new_n2296_;
  assign new_n2612_ = new_n2296_;
  assign new_n2613_ = ~new_n2299_;
  assign new_n2614_ = ~new_n2011_ | ~new_n2312_;
  assign new_n2615_ = ~new_n2302_;
  assign new_n2616_ = ~new_n2305_;
  assign new_n2617_ = ~new_n2306_;
  assign new_n2618_ = new_n2301_ & new_n1462_;
  assign new_n2619_ = ~new_n2308_;
  assign new_n2620_ = ~new_n2035_ | ~new_n2309_;
  assign new_n2621_ = ~new_n2038_ | ~new_n2311_;
  assign new_n2622_ = new_n2303_ & new_n1479_ & new_n2304_ & new_n2301_;
  assign new_n2623_ = ~new_n2040_ | ~new_n2300_;
  assign new_n2624_ = ~new_n2313_;
  assign new_n2625_ = new_n1488_ & new_n2303_ & new_n2301_;
  assign new_n2626_ = ~new_n2314_;
  assign new_n2627_ = new_n2295_ & new_n1494_ & new_n2294_ & new_n2279_;
  assign new_n2628_ = new_n1501_ & new_n2295_ & new_n2279_;
  assign new_n2629_ = new_n2279_ & new_n1506_;
  assign new_n2630_ = new_n2295_ & new_n1509_ & new_n2279_ & new_n2297_ & new_n2294_;
  assign new_n2631_ = new_n2101_ & new_n1830_ & new_n2105_ & new_n2102_;
  assign new_n2632_ = new_n2101_ & new_n1830_ & new_n2098_ & new_n2105_ & new_n2102_;
  assign new_n2633_ = new_n2105_ & new_n1830_;
  assign new_n2634_ = new_n1830_ & new_n2105_ & new_n2102_;
  assign new_n2635_ = new_n2100_ & new_n1831_ & new_n2104_ & new_n2103_;
  assign new_n2636_ = new_n2100_ & new_n1831_ & new_n2099_ & new_n2104_ & new_n2103_;
  assign new_n2637_ = new_n2100_ & new_n1831_ & new_n2104_ & new_n2103_;
  assign new_n2638_ = new_n1831_ & new_n2104_ & new_n2103_;
  assign new_n2639_ = new_n2104_ & new_n1831_;
  assign new_n2640_ = new_n1831_ & new_n2104_ & new_n2103_;
  assign new_n2641_ = ~new_n2054_ | ~new_n2318_;
  assign new_n2642_ = ~new_n2056_ | ~new_n2319_;
  assign new_n2643_ = new_n2322_ & new_n2061_ & new_n2059_;
  assign new_n2644_ = new_n2321_ & new_n2323_ & new_n2320_;
  assign new_n2645_ = ~new_n2321_;
  assign new_n2646_ = ~new_n2322_;
  assign new_n2647_ = ~new_n2063_ | ~new_n2325_;
  assign new_n2648_ = ~new_n2064_ | ~new_n2324_;
  assign new_n2649_ = ~new_n2065_ | ~new_n2327_;
  assign new_n2650_ = ~new_n2066_ | ~new_n2326_;
  assign new_n2651_ = new_n2328_ & new_n2330_ & new_n2331_;
  assign new_n2652_ = ~new_n2328_;
  assign new_n2653_ = ~new_n2329_;
  assign new_n2654_ = new_n2329_ & new_n2068_ & new_n2069_;
  assign new_n2655_ = new_n1571_ & new_n2544_;
  assign new_n2656_ = pi205 & new_n2641_;
  assign new_n2657_ = new_n2105_ & pi205 & new_n2641_;
  assign new_n2658_ = new_n2105_ & new_n2102_ & pi205 & new_n2641_;
  assign new_n2659_ = new_n2101_ & new_n2105_ & new_n2102_ & pi205 & new_n2641_;
  assign new_n2660_ = new_n2359_ | new_n2347_ | new_n1216_ | new_n2339_;
  assign new_n2661_ = new_n2365_ | new_n2351_ | new_n1217_ | new_n2340_;
  assign new_n2662_ = new_n2333_ & new_n2373_;
  assign new_n2663_ = ~new_n2334_;
  assign new_n2664_ = ~new_n2335_;
  assign new_n2665_ = ~new_n2336_;
  assign new_n2666_ = ~new_n2337_;
  assign new_n2667_ = new_n2338_ & new_n2374_;
  assign new_n2668_ = ~new_n2360_ & ~new_n1218_ & ~new_n2349_;
  assign new_n2669_ = new_n2343_ | new_n2361_ | new_n1218_ | new_n2348_;
  assign new_n2670_ = ~new_n2366_ & ~new_n1219_ & ~new_n2350_;
  assign new_n2671_ = new_n2345_ | new_n2364_ | new_n1219_ | new_n2352_;
  assign new_n2672_ = ~new_n2341_;
  assign new_n2673_ = ~new_n2342_;
  assign new_n2674_ = ~new_n2344_;
  assign new_n2675_ = ~new_n2346_;
  assign new_n2676_ = ~new_n1220_ & ~new_n2363_;
  assign new_n2677_ = new_n2355_ | new_n1220_ | new_n2362_;
  assign new_n2678_ = new_n1221_ | new_n2367_;
  assign new_n2679_ = ~new_n2353_;
  assign new_n2680_ = ~new_n2354_;
  assign new_n2681_ = ~new_n2357_;
  assign new_n2682_ = ~new_n2358_;
  assign new_n2683_ = ~new_n2353_ | ~new_n1877_;
  assign new_n2684_ = ~new_n2368_;
  assign new_n2685_ = ~new_n2369_;
  assign new_n2686_ = ~new_n2354_ | ~new_n1583_;
  assign new_n2687_ = new_n2404_ | new_n2392_ | new_n2383_ | new_n1226_ | new_n2376_;
  assign new_n2688_ = new_n2408_ | new_n2396_ | new_n2386_ | new_n1227_ | new_n2377_;
  assign new_n2689_ = ~new_n2371_;
  assign new_n2690_ = ~new_n2372_;
  assign new_n2691_ = ~new_n2373_;
  assign new_n2692_ = ~new_n2375_;
  assign new_n2693_ = ~new_n2409_ & ~new_n2394_ & ~new_n1229_ & ~new_n2384_;
  assign new_n2694_ = new_n2380_ | new_n2407_ | new_n2395_ | new_n1229_ | new_n2385_;
  assign new_n2695_ = ~new_n2378_;
  assign new_n2696_ = ~new_n2379_;
  assign new_n2697_ = ~new_n2381_;
  assign new_n2698_ = ~new_n2412_ & ~new_n1231_ & ~new_n2397_;
  assign new_n2699_ = new_n2389_ | new_n2410_ | new_n1231_ | new_n2398_;
  assign new_n2700_ = ~new_n2387_;
  assign new_n2701_ = ~new_n2388_;
  assign new_n2702_ = ~new_n2390_;
  assign new_n2703_ = new_n1233_ | new_n2411_;
  assign new_n2704_ = ~new_n2399_;
  assign new_n2705_ = ~new_n2400_;
  assign new_n2706_ = ~new_n2402_;
  assign new_n2707_ = ~new_n2413_;
  assign new_n2708_ = ~new_n2414_;
  assign new_n2709_ = ~new_n2415_;
  assign new_n2710_ = new_n2442_ | new_n2430_ | new_n1237_ | new_n2422_;
  assign new_n2711_ = new_n2448_ | new_n2434_ | new_n1238_ | new_n2423_;
  assign new_n2712_ = ~new_n2416_;
  assign new_n2713_ = ~new_n2417_;
  assign new_n2714_ = ~new_n2418_;
  assign new_n2715_ = ~new_n2419_;
  assign new_n2716_ = ~new_n2420_;
  assign new_n2717_ = ~new_n2421_;
  assign new_n2718_ = ~new_n2443_ & ~new_n1239_ & ~new_n2432_;
  assign new_n2719_ = new_n2426_ | new_n2444_ | new_n1239_ | new_n2431_;
  assign new_n2720_ = ~new_n2449_ & ~new_n1240_ & ~new_n2433_;
  assign new_n2721_ = new_n2428_ | new_n2447_ | new_n1240_ | new_n2435_;
  assign new_n2722_ = ~new_n2424_;
  assign new_n2723_ = ~new_n2425_;
  assign new_n2724_ = ~new_n2427_;
  assign new_n2725_ = ~new_n2429_;
  assign new_n2726_ = ~new_n1241_ & ~new_n2446_;
  assign new_n2727_ = new_n2441_ | new_n1241_ | new_n2445_;
  assign new_n2728_ = new_n1242_ | new_n2450_;
  assign new_n2729_ = ~new_n2437_;
  assign new_n2730_ = ~new_n2438_;
  assign new_n2731_ = ~new_n2439_;
  assign new_n2732_ = ~new_n2440_;
  assign new_n2733_ = ~new_n2439_ | ~new_n1898_;
  assign new_n2734_ = ~new_n2451_;
  assign new_n2735_ = ~new_n2452_;
  assign new_n2736_ = ~new_n2440_ | ~new_n1607_;
  assign new_n2737_ = new_n2632_ | new_n2471_ | new_n2463_ | new_n1247_ | new_n2457_;
  assign new_n2738_ = new_n2636_ | new_n2475_ | new_n2466_ | new_n1248_ | new_n2458_;
  assign new_n2739_ = new_n2105_ & new_n2098_ & new_n2102_ & new_n2101_ & new_n2641_;
  assign new_n2740_ = ~new_n2454_;
  assign new_n2741_ = ~new_n2455_;
  assign new_n2742_ = ~new_n2456_;
  assign new_n2743_ = new_n2099_ & new_n2100_ & new_n2103_ & new_n2642_ & new_n2104_;
  assign new_n2744_ = ~new_n2637_ & ~new_n2473_ & ~new_n1250_ & ~new_n2464_;
  assign new_n2745_ = ~new_n2459_;
  assign new_n2746_ = new_n2104_ & new_n2100_ & new_n2642_ & new_n2103_;
  assign new_n2747_ = ~new_n2460_;
  assign new_n2748_ = ~new_n2461_;
  assign new_n2749_ = ~new_n2640_ & ~new_n1252_ & ~new_n2476_;
  assign new_n2750_ = ~new_n2467_;
  assign new_n2751_ = ~new_n2468_;
  assign new_n2752_ = ~new_n2469_;
  assign new_n2753_ = new_n2104_ & new_n2642_ & new_n2103_;
  assign new_n2754_ = new_n1254_ | new_n2639_;
  assign new_n2755_ = ~new_n2478_;
  assign new_n2756_ = ~new_n2479_;
  assign new_n2757_ = new_n2642_ & new_n2104_;
  assign new_n2758_ = ~new_n2480_;
  assign new_n2759_ = ~new_n2503_ | ~new_n2482_;
  assign new_n2760_ = new_n2107_ & new_n2512_;
  assign new_n2761_ = new_n2108_ & new_n2516_;
  assign new_n2762_ = ~new_n2493_ | ~new_n2489_;
  assign new_n2763_ = ~new_n2492_ | ~new_n2490_;
  assign new_n2764_ = new_n2520_ & new_n2113_;
  assign new_n2765_ = ~new_n2492_;
  assign new_n2766_ = ~new_n2493_;
  assign new_n2767_ = ~new_n2501_ | ~new_n2494_;
  assign new_n2768_ = ~new_n2502_ | ~new_n2495_;
  assign new_n2769_ = ~new_n2496_;
  assign new_n2770_ = ~new_n2497_;
  assign new_n2771_ = ~new_n2500_;
  assign new_n2772_ = ~new_n2501_;
  assign new_n2773_ = ~new_n2502_;
  assign new_n2774_ = new_n2500_ | new_n2131_;
  assign new_n2775_ = ~new_n1268_ | ~new_n2506_;
  assign new_n2776_ = ~new_n993_ | ~new_n2507_;
  assign new_n2777_ = ~new_n2516_;
  assign new_n2778_ = ~new_n2522_;
  assign new_n2779_ = ~new_n2523_;
  assign new_n2780_ = ~new_n2527_;
  assign new_n2781_ = ~new_n2528_;
  assign new_n2782_ = new_n2515_ & new_n2202_ & new_n1931_;
  assign new_n2783_ = ~new_n2533_;
  assign new_n2784_ = new_n2533_ | new_n2187_;
  assign new_n2785_ = ~new_n2527_ | ~new_n1650_;
  assign new_n2786_ = ~new_n2528_ | ~new_n1292_;
  assign new_n2787_ = new_n2514_ & new_n1939_ & new_n2171_;
  assign new_n2788_ = ~new_n2620_ | ~new_n1658_;
  assign new_n2789_ = ~new_n2621_ | ~new_n1946_;
  assign new_n2790_ = new_n2543_ & new_n1305_;
  assign new_n2791_ = new_n1308_ & new_n2542_;
  assign new_n2792_ = ~new_n2542_;
  assign new_n2793_ = ~new_n2544_;
  assign new_n2794_ = ~new_n2552_;
  assign new_n2795_ = ~new_n2553_;
  assign new_n2796_ = ~new_n2557_;
  assign new_n2797_ = new_n2547_ & new_n2247_ & new_n1957_;
  assign new_n2798_ = new_n2557_ | new_n2233_;
  assign new_n2799_ = ~new_n2590_ | ~new_n1678_;
  assign new_n2800_ = ~new_n2591_ | ~new_n1328_;
  assign new_n2801_ = new_n2546_ & new_n1960_ & new_n2229_;
  assign new_n2802_ = new_n2568_ & new_n1963_ & new_n2250_;
  assign new_n2803_ = new_n2567_ & new_n2249_ & new_n1964_;
  assign new_n2804_ = new_n2572_ & new_n1966_ & new_n2254_;
  assign new_n2805_ = new_n2571_ & new_n2253_ & new_n1967_;
  assign new_n2806_ = ~new_n2257_ | ~new_n2580_;
  assign new_n2807_ = new_n2575_ & new_n2595_;
  assign new_n2808_ = ~new_n2575_;
  assign new_n2809_ = ~new_n2259_ | ~new_n2578_;
  assign new_n2810_ = ~new_n2261_ | ~new_n2576_;
  assign new_n2811_ = ~new_n2263_ | ~new_n2573_;
  assign new_n2812_ = new_n2581_ & new_n2600_ & new_n2589_;
  assign new_n2813_ = ~new_n2581_;
  assign new_n2814_ = ~new_n2582_;
  assign new_n2815_ = new_n2606_ & new_n2584_;
  assign new_n2816_ = new_n2585_ & new_n2602_ & new_n2588_;
  assign new_n2817_ = ~new_n2585_;
  assign new_n2818_ = ~new_n2586_;
  assign new_n2819_ = new_n2586_ & new_n2285_ & new_n2268_;
  assign new_n2820_ = new_n2582_ & new_n2283_ & new_n2269_;
  assign new_n2821_ = ~new_n2590_;
  assign new_n2822_ = ~new_n2591_;
  assign new_n2823_ = new_n2630_ | new_n2627_ | new_n2628_ | new_n1393_ | new_n2629_;
  assign new_n2824_ = ~new_n2596_;
  assign new_n2825_ = ~new_n2597_;
  assign new_n2826_ = ~new_n2598_;
  assign new_n2827_ = new_n2599_ & new_n2626_ & new_n2619_;
  assign new_n2828_ = ~new_n2599_;
  assign new_n2829_ = new_n2574_ | new_n2577_ | new_n1402_ | new_n2579_;
  assign new_n2830_ = ~new_n2595_ | ~pi048;
  assign new_n2831_ = ~new_n2604_;
  assign new_n2832_ = new_n2605_ & new_n2608_ & new_n2609_;
  assign new_n2833_ = ~new_n2605_;
  assign new_n2834_ = ~new_n2606_;
  assign new_n2835_ = ~new_n2290_ | ~new_n2615_;
  assign new_n2836_ = new_n2604_ & new_n2291_ & new_n2292_;
  assign new_n2837_ = ~new_n2611_;
  assign new_n2838_ = ~new_n2612_;
  assign new_n2839_ = new_n2612_ & new_n2293_ & new_n2009_;
  assign new_n2840_ = new_n2611_ & new_n2610_ & new_n2298_;
  assign new_n2841_ = ~new_n2299_ | ~new_n2624_;
  assign new_n2842_ = new_n2622_ | new_n2625_ | new_n1439_ | new_n2618_;
  assign new_n2843_ = ~new_n2623_ | ~new_n2614_;
  assign new_n2844_ = ~new_n2302_ | ~new_n2607_;
  assign new_n2845_ = ~new_n2305_ | ~new_n2617_;
  assign new_n2846_ = ~new_n2306_ | ~new_n2616_;
  assign new_n2847_ = new_n2587_ | new_n2601_ | new_n2603_ | new_n1465_ | new_n2583_;
  assign new_n2848_ = new_n2597_ & new_n2046_ & new_n2032_;
  assign new_n2849_ = new_n2596_ & new_n2315_ & new_n2307_;
  assign new_n2850_ = new_n2598_ & new_n2314_ & new_n2308_;
  assign new_n2851_ = ~new_n2620_;
  assign new_n2852_ = ~new_n2621_;
  assign new_n2853_ = ~new_n2313_ | ~new_n2613_;
  assign new_n2854_ = new_n2641_;
  assign new_n2855_ = new_n2642_;
  assign new_n2856_ = new_n2642_;
  assign new_n2857_ = new_n2645_ & new_n2059_ & new_n2323_;
  assign new_n2858_ = new_n2646_ & new_n2320_ & new_n2061_;
  assign new_n2859_ = ~new_n2648_ | ~new_n2647_;
  assign new_n2860_ = ~new_n2649_ | ~new_n2650_;
  assign new_n2861_ = new_n2653_ & new_n2331_ & new_n2068_;
  assign new_n2862_ = new_n2652_ & new_n2069_ & new_n2330_;
  assign new_n2863_ = ~new_n2854_ | ~new_n425_;
  assign new_n2864_ = ~new_n2743_ | ~pi205;
  assign new_n2865_ = new_n2739_ & pi205;
  assign new_n2866_ = new_n2333_ & new_n2688_;
  assign new_n2867_ = ~new_n2669_ | ~new_n2665_;
  assign new_n2868_ = ~new_n2668_ | ~new_n2666_;
  assign new_n2869_ = new_n2687_ & new_n2338_;
  assign new_n2870_ = ~new_n2668_;
  assign new_n2871_ = ~new_n2669_;
  assign new_n2872_ = ~new_n2670_;
  assign new_n2873_ = ~new_n2671_;
  assign new_n2874_ = ~new_n2676_ | ~new_n2672_;
  assign new_n2875_ = ~new_n2677_ | ~new_n2673_;
  assign new_n2876_ = ~new_n2676_;
  assign new_n2877_ = ~new_n2677_;
  assign new_n2878_ = ~new_n2678_;
  assign new_n2879_ = new_n2678_ | new_n2356_;
  assign new_n2880_ = ~new_n1578_ | ~new_n2679_;
  assign new_n2881_ = ~new_n1225_ | ~new_n2680_;
  assign new_n2882_ = ~new_n2688_;
  assign new_n2883_ = ~new_n2693_;
  assign new_n2884_ = ~new_n2694_;
  assign new_n2885_ = ~new_n2698_;
  assign new_n2886_ = ~new_n2699_;
  assign new_n2887_ = ~new_n2703_;
  assign new_n2888_ = new_n2703_ | new_n2401_;
  assign new_n2889_ = ~new_n2698_ | ~new_n1889_;
  assign new_n2890_ = ~new_n2699_ | ~new_n1594_;
  assign new_n2891_ = ~new_n2710_;
  assign new_n2892_ = ~new_n2711_;
  assign new_n2893_ = new_n2416_ & new_n2738_;
  assign new_n2894_ = new_n2416_ & new_n2743_;
  assign new_n2895_ = ~new_n2719_ | ~new_n2715_;
  assign new_n2896_ = ~new_n2718_ | ~new_n2716_;
  assign new_n2897_ = new_n2421_ & new_n2739_;
  assign new_n2898_ = new_n2737_ & new_n2421_;
  assign new_n2899_ = ~new_n2718_;
  assign new_n2900_ = ~new_n2719_;
  assign new_n2901_ = ~new_n2720_;
  assign new_n2902_ = ~new_n2721_;
  assign new_n2903_ = ~new_n2726_ | ~new_n2722_;
  assign new_n2904_ = ~new_n2727_ | ~new_n2723_;
  assign new_n2905_ = ~new_n2726_;
  assign new_n2906_ = ~new_n2727_;
  assign new_n2907_ = ~new_n2728_;
  assign new_n2908_ = new_n2728_ | new_n2436_;
  assign new_n2909_ = ~new_n1602_ | ~new_n2731_;
  assign new_n2910_ = ~new_n1246_ | ~new_n2732_;
  assign new_n2911_ = ~new_n2738_;
  assign new_n2912_ = ~new_n2743_;
  assign new_n2913_ = new_n2659_ | new_n2631_ | new_n2470_ | new_n1249_ | new_n2462_;
  assign new_n2914_ = ~new_n2744_;
  assign new_n2915_ = new_n2746_ | new_n2635_ | new_n2474_ | new_n1250_ | new_n2465_;
  assign new_n2916_ = new_n2658_ | new_n2634_ | new_n1251_ | new_n2472_;
  assign new_n2917_ = ~new_n2749_;
  assign new_n2918_ = new_n2753_ | new_n2638_ | new_n1252_ | new_n2477_;
  assign new_n2919_ = new_n2657_ | new_n1253_ | new_n2633_;
  assign new_n2920_ = new_n2754_ | new_n2757_;
  assign new_n2921_ = ~new_n2754_;
  assign new_n2922_ = new_n2481_ | new_n2760_;
  assign new_n2923_ = ~new_n2759_;
  assign new_n2924_ = new_n2487_ | new_n2761_;
  assign new_n2925_ = new_n2488_ | new_n2764_;
  assign new_n2926_ = ~new_n2111_ | ~new_n2766_;
  assign new_n2927_ = ~new_n2112_ | ~new_n2765_;
  assign new_n2928_ = ~new_n2116_ | ~new_n2772_;
  assign new_n2929_ = ~new_n2117_ | ~new_n2773_;
  assign new_n2930_ = ~new_n2771_;
  assign new_n2931_ = ~new_n2774_;
  assign new_n2932_ = ~new_n2771_ | ~new_n1628_;
  assign new_n2933_ = ~new_n2508_ | ~new_n2775_;
  assign new_n2934_ = ~new_n2509_ | ~new_n2776_;
  assign new_n2935_ = ~new_n2774_ | ~new_n1271_;
  assign new_n2936_ = ~new_n2787_ & ~new_n2513_;
  assign new_n2937_ = new_n2777_ & new_n2519_;
  assign new_n2938_ = ~new_n2782_ & ~new_n2529_;
  assign new_n2939_ = ~new_n2783_;
  assign new_n2940_ = ~new_n2784_;
  assign new_n2941_ = ~new_n1291_ | ~new_n2780_;
  assign new_n2942_ = ~new_n1020_ | ~new_n2781_;
  assign new_n2943_ = ~new_n1300_ | ~new_n2851_;
  assign new_n2944_ = new_n1301_ | new_n2791_;
  assign new_n2945_ = ~new_n1660_ | ~new_n2852_;
  assign new_n2946_ = new_n1302_ | new_n2790_;
  assign new_n2947_ = ~new_n2801_ & ~new_n2545_;
  assign new_n2948_ = new_n2792_ & new_n2550_;
  assign new_n2949_ = ~new_n2796_;
  assign new_n2950_ = ~new_n2797_ & ~new_n2559_;
  assign new_n2951_ = ~new_n2798_;
  assign new_n2952_ = ~new_n1327_ | ~new_n2821_;
  assign new_n2953_ = ~new_n1050_ | ~new_n2822_;
  assign new_n2954_ = ~new_n2803_ & ~new_n2565_;
  assign new_n2955_ = ~new_n2802_ & ~new_n2566_;
  assign new_n2956_ = ~new_n2805_ & ~new_n2569_;
  assign new_n2957_ = ~new_n2804_ & ~new_n2570_;
  assign new_n2958_ = ~new_n2806_ | ~new_n2811_;
  assign new_n2959_ = new_n2575_ & new_n2823_;
  assign new_n2960_ = ~new_n2809_ | ~new_n2810_;
  assign new_n2961_ = new_n2817_ & new_n2268_ & new_n2602_;
  assign new_n2962_ = new_n2813_ & new_n2269_ & new_n2600_;
  assign new_n2963_ = ~new_n2823_;
  assign new_n2964_ = ~new_n2829_;
  assign new_n2965_ = new_n2814_ & new_n2589_ & new_n2283_;
  assign new_n2966_ = new_n2818_ & new_n2588_ & new_n2285_;
  assign new_n2967_ = new_n2332_ & new_n2483_ & new_n2815_ & pi048 & new_n2807_;
  assign new_n2968_ = new_n2483_ & new_n2815_ & pi048 & new_n2807_;
  assign new_n2969_ = new_n2332_ & new_n2483_ & new_n2815_ & pi048 & new_n2807_;
  assign new_n2970_ = new_n2606_ & new_n2847_;
  assign new_n2971_ = ~new_n2835_ | ~new_n2844_;
  assign new_n2972_ = new_n2831_ & new_n2609_ & new_n2291_;
  assign new_n2973_ = new_n2833_ & new_n2292_ & new_n2608_;
  assign new_n2974_ = new_n2838_ & new_n2298_ & new_n2293_;
  assign new_n2975_ = new_n2837_ & new_n2009_ & new_n2610_;
  assign new_n2976_ = ~new_n2853_ | ~new_n2841_;
  assign new_n2977_ = ~new_n2842_;
  assign new_n2978_ = ~new_n2843_;
  assign new_n2979_ = ~new_n2846_ | ~new_n2845_;
  assign new_n2980_ = ~new_n2847_;
  assign new_n2981_ = new_n2824_ & new_n2032_ & new_n2315_;
  assign new_n2982_ = new_n2828_ & new_n2308_ & new_n2626_;
  assign new_n2983_ = new_n1807_ | new_n2655_;
  assign new_n2984_ = new_n2826_ & new_n2619_ & new_n2314_;
  assign new_n2985_ = new_n2825_ & new_n2307_ & new_n2046_;
  assign new_n2986_ = new_n1830_ | new_n2656_;
  assign new_n2987_ = ~new_n2749_ | ~new_n2317_;
  assign new_n2988_ = ~new_n2854_;
  assign new_n2989_ = ~new_n2855_;
  assign new_n2990_ = ~new_n2856_;
  assign new_n2991_ = ~new_n2858_ & ~new_n2643_;
  assign new_n2992_ = ~new_n2857_ & ~new_n2644_;
  assign new_n2993_ = ~new_n2859_;
  assign new_n2994_ = ~new_n2860_;
  assign new_n2995_ = ~new_n2862_ & ~new_n2651_;
  assign new_n2996_ = ~new_n2861_ & ~new_n2654_;
  assign new_n2997_ = new_n2922_ & new_n2332_;
  assign new_n2998_ = new_n2922_ & new_n2332_;
  assign new_n2999_ = ~new_n316_ | ~new_n2988_;
  assign new_n3000_ = new_n2667_ & pi205 & new_n2897_;
  assign new_n3001_ = new_n2491_ & new_n2667_ & pi205 & new_n2897_;
  assign new_n3002_ = new_n2911_ & new_n2864_;
  assign new_n3003_ = new_n2662_ & pi205 & new_n2894_;
  assign new_n3004_ = new_n2484_ & new_n2662_ & pi205 & new_n2894_;
  assign new_n3005_ = new_n2541_ & new_n2484_ & new_n2662_ & pi205 & new_n2894_;
  assign new_n3006_ = new_n2540_ & new_n2491_ & new_n2667_ & pi205 & new_n2897_;
  assign new_n3007_ = new_n2660_ | new_n2869_;
  assign new_n3008_ = new_n2661_ | new_n2866_;
  assign new_n3009_ = ~new_n2336_ | ~new_n2871_;
  assign new_n3010_ = ~new_n2337_ | ~new_n2870_;
  assign new_n3011_ = ~new_n2341_ | ~new_n2876_;
  assign new_n3012_ = ~new_n2342_ | ~new_n2877_;
  assign new_n3013_ = ~new_n2878_;
  assign new_n3014_ = ~new_n2879_;
  assign new_n3015_ = ~new_n2683_ | ~new_n2880_;
  assign new_n3016_ = ~new_n2878_ | ~new_n1878_;
  assign new_n3017_ = ~new_n2879_ | ~new_n1580_;
  assign new_n3018_ = ~new_n2686_ | ~new_n2881_;
  assign new_n3019_ = new_n2882_ & new_n2691_;
  assign new_n3020_ = ~new_n2887_;
  assign new_n3021_ = ~new_n2888_;
  assign new_n3022_ = ~new_n1592_ | ~new_n2885_;
  assign new_n3023_ = ~new_n1236_ | ~new_n2886_;
  assign new_n3024_ = new_n2710_ | new_n2898_;
  assign new_n3025_ = new_n2711_ | new_n2893_;
  assign new_n3026_ = ~new_n2892_ | ~new_n2712_;
  assign new_n3027_ = ~new_n2419_ | ~new_n2900_;
  assign new_n3028_ = ~new_n2420_ | ~new_n2899_;
  assign new_n3029_ = ~new_n2891_ | ~new_n2717_;
  assign new_n3030_ = ~new_n2424_ | ~new_n2905_;
  assign new_n3031_ = ~new_n2425_ | ~new_n2906_;
  assign new_n3032_ = ~new_n2907_;
  assign new_n3033_ = ~new_n2908_;
  assign new_n3034_ = ~new_n2733_ | ~new_n2909_;
  assign new_n3035_ = ~new_n2907_ | ~new_n1899_;
  assign new_n3036_ = ~new_n2908_ | ~new_n1604_;
  assign new_n3037_ = ~new_n2736_ | ~new_n2910_;
  assign new_n3038_ = new_n2737_ | new_n2865_;
  assign new_n3039_ = new_n2911_ & new_n2912_;
  assign new_n3040_ = ~new_n2913_ | ~new_n2740_;
  assign new_n3041_ = ~new_n2913_;
  assign new_n3042_ = ~new_n2915_;
  assign new_n3043_ = ~new_n2916_ | ~new_n2748_;
  assign new_n3044_ = ~new_n2916_;
  assign new_n3045_ = ~new_n2918_;
  assign new_n3046_ = ~new_n2919_ | ~new_n2750_;
  assign new_n3047_ = ~new_n2919_;
  assign new_n3048_ = ~new_n2920_;
  assign new_n3049_ = ~new_n2921_;
  assign new_n3050_ = ~new_n2986_ | ~new_n2758_;
  assign new_n3051_ = ~new_n2926_ | ~new_n2762_;
  assign new_n3052_ = ~new_n2927_ | ~new_n2763_;
  assign new_n3053_ = ~new_n2928_ | ~new_n2767_;
  assign new_n3054_ = ~new_n2929_ | ~new_n2768_;
  assign new_n3055_ = ~new_n1267_ | ~new_n2930_;
  assign new_n3056_ = ~new_n2934_;
  assign new_n3057_ = ~new_n994_ | ~new_n2931_;
  assign new_n3058_ = ~new_n2936_ | ~new_n2938_;
  assign new_n3059_ = ~new_n2937_;
  assign new_n3060_ = ~new_n2785_ | ~new_n2941_;
  assign new_n3061_ = ~new_n2786_ | ~new_n2942_;
  assign new_n3062_ = ~new_n2943_ | ~new_n2788_;
  assign new_n3063_ = ~new_n2945_ | ~new_n2789_;
  assign new_n3064_ = new_n2925_ & new_n2540_;
  assign new_n3065_ = new_n2924_ & new_n2541_;
  assign new_n3066_ = ~new_n2947_ | ~new_n2950_;
  assign new_n3067_ = ~new_n2948_;
  assign new_n3068_ = ~new_n2799_ | ~new_n2952_;
  assign new_n3069_ = ~new_n2800_ | ~new_n2953_;
  assign new_n3070_ = ~new_n2955_ | ~new_n2954_;
  assign new_n3071_ = ~new_n2957_ | ~new_n2956_;
  assign new_n3072_ = ~new_n2958_;
  assign new_n3073_ = ~new_n2964_ | ~new_n2808_;
  assign new_n3074_ = ~new_n2960_;
  assign new_n3075_ = ~new_n2962_ & ~new_n2812_;
  assign new_n3076_ = ~new_n2961_ & ~new_n2816_;
  assign new_n3077_ = ~new_n2966_ & ~new_n2819_;
  assign new_n3078_ = ~new_n2965_ & ~new_n2820_;
  assign new_n3079_ = ~new_n2982_ & ~new_n2827_;
  assign new_n3080_ = new_n2829_ | new_n2959_;
  assign new_n3081_ = new_n2963_ & new_n2830_;
  assign new_n3082_ = ~new_n2973_ & ~new_n2832_;
  assign new_n3083_ = ~new_n2977_ | ~new_n2834_;
  assign new_n3084_ = ~new_n2971_;
  assign new_n3085_ = ~new_n2972_ & ~new_n2836_;
  assign new_n3086_ = ~new_n2974_ & ~new_n2839_;
  assign new_n3087_ = ~new_n2975_ & ~new_n2840_;
  assign new_n3088_ = ~new_n2976_;
  assign new_n3089_ = new_n2842_ | new_n2970_;
  assign new_n3090_ = ~new_n2979_;
  assign new_n3091_ = ~new_n2985_ & ~new_n2848_;
  assign new_n3092_ = ~new_n2981_ & ~new_n2849_;
  assign new_n3093_ = ~new_n2984_ & ~new_n2850_;
  assign new_n3094_ = ~new_n2986_;
  assign new_n3095_ = ~new_n2053_ | ~new_n2917_;
  assign new_n3096_ = ~new_n2918_ | ~new_n2055_;
  assign new_n3097_ = ~new_n2992_ | ~new_n2991_;
  assign new_n3098_ = ~new_n2995_ | ~new_n2996_;
  assign new_n3099_ = new_n2332_ & new_n3089_ & new_n2483_;
  assign new_n3100_ = new_n2332_ & new_n2483_ & new_n3080_ & new_n2815_;
  assign new_n3101_ = new_n2332_ & new_n3089_ & new_n2483_;
  assign new_n3102_ = new_n2332_ & new_n2483_ & new_n3080_ & new_n2815_;
  assign po056 = ~new_n2863_ | ~new_n2999_;
  assign new_n3104_ = ~new_n3002_;
  assign new_n3105_ = new_n3025_ & new_n2662_;
  assign new_n3106_ = ~new_n3009_ | ~new_n2867_;
  assign new_n3107_ = ~new_n3010_ | ~new_n2868_;
  assign new_n3108_ = new_n3024_ & new_n2667_;
  assign new_n3109_ = ~new_n3011_ | ~new_n2874_;
  assign new_n3110_ = ~new_n3012_ | ~new_n2875_;
  assign new_n3111_ = ~new_n1579_ | ~new_n3013_;
  assign new_n3112_ = ~new_n1224_ | ~new_n3014_;
  assign new_n3113_ = ~new_n3018_;
  assign new_n3114_ = ~new_n3019_;
  assign new_n3115_ = ~new_n2889_ | ~new_n3022_;
  assign new_n3116_ = ~new_n2890_ | ~new_n3023_;
  assign new_n3117_ = new_n3002_ & new_n2711_;
  assign new_n3118_ = ~new_n3027_ | ~new_n2895_;
  assign new_n3119_ = ~new_n3028_ | ~new_n2896_;
  assign new_n3120_ = new_n3029_ & new_n3038_;
  assign new_n3121_ = ~new_n3030_ | ~new_n2903_;
  assign new_n3122_ = ~new_n3031_ | ~new_n2904_;
  assign new_n3123_ = ~new_n1603_ | ~new_n3032_;
  assign new_n3124_ = ~new_n1245_ | ~new_n3033_;
  assign new_n3125_ = new_n3038_ & new_n2453_;
  assign new_n3126_ = ~new_n3037_;
  assign new_n3127_ = ~new_n3038_;
  assign new_n3128_ = ~new_n3039_;
  assign new_n3129_ = ~new_n2454_ | ~new_n3041_;
  assign new_n3130_ = ~new_n2461_ | ~new_n3044_;
  assign new_n3131_ = ~new_n2467_ | ~new_n3047_;
  assign new_n3132_ = ~new_n2480_ | ~new_n3094_;
  assign new_n3133_ = ~new_n3058_ | ~new_n2923_;
  assign new_n3134_ = new_n3089_ & new_n2483_;
  assign new_n3135_ = new_n2483_ & new_n3080_ & new_n2815_;
  assign new_n3136_ = new_n2541_ & new_n3008_ & new_n2484_;
  assign new_n3137_ = new_n2541_ & new_n2484_ & new_n3025_ & new_n2662_;
  assign new_n3138_ = new_n3008_ & new_n2484_;
  assign new_n3139_ = new_n2484_ & new_n3025_ & new_n2662_;
  assign new_n3140_ = ~new_n3052_;
  assign new_n3141_ = new_n2540_ & new_n3007_ & new_n2491_;
  assign new_n3142_ = new_n2540_ & new_n2491_ & new_n3024_ & new_n2667_;
  assign new_n3143_ = new_n3007_ & new_n2491_;
  assign new_n3144_ = new_n2491_ & new_n3024_ & new_n2667_;
  assign new_n3145_ = ~new_n3053_;
  assign new_n3146_ = ~new_n2932_ | ~new_n3055_;
  assign new_n3147_ = ~new_n2935_ | ~new_n3057_;
  assign new_n3148_ = ~new_n3058_;
  assign new_n3149_ = ~new_n3060_ | ~new_n2939_;
  assign new_n3150_ = ~new_n3061_ | ~new_n2940_;
  assign new_n3151_ = ~new_n3060_;
  assign new_n3152_ = ~new_n3061_;
  assign new_n3153_ = ~new_n3066_ | ~new_n1942_;
  assign new_n3154_ = ~new_n3062_;
  assign new_n3155_ = ~new_n3063_;
  assign new_n3156_ = ~new_n3062_ | ~new_n1664_;
  assign new_n3157_ = ~new_n3063_ | ~new_n1665_;
  assign new_n3158_ = ~new_n3066_;
  assign new_n3159_ = ~new_n3068_ | ~new_n2949_;
  assign new_n3160_ = ~new_n3069_ | ~new_n2951_;
  assign new_n3161_ = ~new_n3068_;
  assign new_n3162_ = ~new_n3069_;
  assign new_n3163_ = ~new_n3070_;
  assign new_n3164_ = ~new_n3071_;
  assign new_n3165_ = ~new_n3075_ | ~new_n3078_;
  assign new_n3166_ = ~new_n3076_ | ~new_n3077_;
  assign new_n3167_ = ~new_n3079_ | ~new_n3093_;
  assign new_n3168_ = new_n3081_ & new_n2829_;
  assign new_n3169_ = ~new_n3081_;
  assign new_n3170_ = ~new_n3082_ | ~new_n3085_;
  assign new_n3171_ = ~new_n3087_ | ~new_n3086_;
  assign new_n3172_ = ~new_n3092_ | ~new_n3091_;
  assign new_n3173_ = ~new_n2987_ | ~new_n3095_;
  assign new_n3174_ = ~new_n1832_ | ~new_n3045_;
  assign new_n3175_ = ~new_n3097_;
  assign new_n3176_ = ~new_n3097_ | ~new_n2062_;
  assign new_n3177_ = ~new_n3070_ | ~new_n2993_;
  assign new_n3178_ = ~new_n3071_ | ~new_n2994_;
  assign new_n3179_ = ~new_n3098_;
  assign new_n3180_ = ~new_n3098_ | ~new_n2070_;
  assign new_n3181_ = new_n3000_ | new_n3007_ | new_n3108_;
  assign new_n3182_ = new_n3003_ | new_n3008_ | new_n3105_;
  assign new_n3183_ = ~new_n3107_;
  assign new_n3184_ = ~new_n3109_;
  assign new_n3185_ = ~new_n3016_ | ~new_n3111_;
  assign new_n3186_ = ~new_n3017_ | ~new_n3112_;
  assign new_n3187_ = ~new_n3115_ | ~new_n3020_;
  assign new_n3188_ = ~new_n3116_ | ~new_n3021_;
  assign new_n3189_ = ~new_n3115_;
  assign new_n3190_ = ~new_n3116_;
  assign new_n3191_ = new_n2710_ & new_n3127_;
  assign new_n3192_ = new_n3026_ & new_n3104_;
  assign new_n3193_ = ~new_n3119_;
  assign new_n3194_ = ~new_n3121_;
  assign new_n3195_ = new_n3034_ & new_n3127_;
  assign new_n3196_ = ~new_n3035_ | ~new_n3123_;
  assign new_n3197_ = ~new_n3036_ | ~new_n3124_;
  assign new_n3198_ = new_n2097_ & new_n3127_;
  assign new_n3199_ = new_n3038_ & new_n3118_;
  assign new_n3200_ = new_n3038_ & new_n3122_;
  assign new_n3201_ = new_n3038_ & new_n3126_;
  assign po061 = ~new_n3129_ | ~new_n3040_;
  assign po062 = ~new_n3130_ | ~new_n3043_;
  assign po063 = ~new_n3131_ | ~new_n3046_;
  assign new_n3205_ = ~new_n3173_ | ~new_n3049_;
  assign po064 = ~new_n3132_ | ~new_n3050_;
  assign new_n3207_ = new_n2968_ | new_n3135_ | new_n2922_ | new_n3134_;
  assign new_n3208_ = ~new_n2759_ | ~new_n3148_;
  assign new_n3209_ = new_n3004_ | new_n3139_ | new_n2924_ | new_n3138_;
  assign new_n3210_ = new_n3001_ | new_n3144_ | new_n2925_ | new_n3143_;
  assign new_n3211_ = ~new_n3146_ | ~new_n2769_;
  assign new_n3212_ = ~new_n3147_ | ~new_n2770_;
  assign new_n3213_ = ~new_n3146_;
  assign new_n3214_ = ~new_n3147_;
  assign new_n3215_ = ~new_n2783_ | ~new_n3151_;
  assign new_n3216_ = ~new_n2784_ | ~new_n3152_;
  assign new_n3217_ = ~new_n1655_ | ~new_n3158_;
  assign po060 = new_n3005_ | new_n3137_ | new_n3136_ | new_n2944_ | new_n3065_;
  assign po057 = new_n3006_ | new_n3142_ | new_n3141_ | new_n2946_ | new_n3064_;
  assign new_n3220_ = ~new_n1312_ | ~new_n3154_;
  assign new_n3221_ = ~new_n1313_ | ~new_n3155_;
  assign new_n3222_ = ~new_n2796_ | ~new_n3161_;
  assign new_n3223_ = ~new_n2798_ | ~new_n3162_;
  assign new_n3224_ = ~new_n3172_ | ~new_n3072_;
  assign new_n3225_ = new_n3073_ & new_n3169_;
  assign new_n3226_ = ~new_n3167_ | ~new_n3074_;
  assign new_n3227_ = ~new_n3165_;
  assign new_n3228_ = ~new_n3166_;
  assign new_n3229_ = ~new_n3167_;
  assign po059 = new_n2967_ | new_n3102_ | new_n3101_ | new_n2983_ | new_n2998_;
  assign po058 = new_n2969_ | new_n3100_ | new_n3099_ | new_n2983_ | new_n2997_;
  assign new_n3232_ = ~new_n3170_;
  assign new_n3233_ = ~new_n3170_ | ~new_n3084_;
  assign new_n3234_ = ~new_n3171_;
  assign new_n3235_ = ~new_n3165_ | ~new_n3088_;
  assign new_n3236_ = ~new_n3166_ | ~new_n2978_;
  assign new_n3237_ = ~new_n3171_ | ~new_n3090_;
  assign new_n3238_ = ~new_n3172_;
  assign new_n3239_ = ~new_n3173_;
  assign new_n3240_ = ~new_n3096_ | ~new_n3174_;
  assign new_n3241_ = ~new_n1845_ | ~new_n3175_;
  assign new_n3242_ = ~new_n2859_ | ~new_n3163_;
  assign new_n3243_ = ~new_n2860_ | ~new_n3164_;
  assign new_n3244_ = ~new_n1868_ | ~new_n3179_;
  assign new_n3245_ = new_n3181_;
  assign new_n3246_ = ~new_n3182_;
  assign new_n3247_ = ~new_n3185_ | ~new_n2872_;
  assign new_n3248_ = ~new_n3186_ | ~new_n2873_;
  assign new_n3249_ = ~new_n3185_;
  assign new_n3250_ = ~new_n3186_;
  assign new_n3251_ = ~new_n2887_ | ~new_n3189_;
  assign new_n3252_ = ~new_n2888_ | ~new_n3190_;
  assign new_n3253_ = new_n3192_ | new_n3117_;
  assign new_n3254_ = new_n3191_ | new_n3120_;
  assign new_n3255_ = ~new_n3196_ | ~new_n2901_;
  assign new_n3256_ = ~new_n3197_ | ~new_n2902_;
  assign po067 = new_n3195_ | new_n3201_;
  assign new_n3258_ = ~new_n3196_;
  assign new_n3259_ = ~new_n3197_;
  assign po068 = new_n3198_ | new_n3125_;
  assign new_n3261_ = new_n3193_ & new_n3127_;
  assign new_n3262_ = new_n3194_ & new_n3127_;
  assign new_n3263_ = ~new_n3240_ | ~new_n3048_;
  assign new_n3264_ = ~new_n2921_ | ~new_n3239_;
  assign new_n3265_ = ~new_n3208_ | ~new_n3133_;
  assign new_n3266_ = new_n3209_;
  assign new_n3267_ = new_n3210_;
  assign new_n3268_ = ~new_n2496_ | ~new_n3213_;
  assign new_n3269_ = ~new_n2497_ | ~new_n3214_;
  assign new_n3270_ = new_n2156_ & new_n3181_;
  assign new_n3271_ = new_n1928_ & new_n1935_ & new_n1934_ & new_n3181_ & new_n1941_;
  assign new_n3272_ = new_n1935_ & new_n1934_ & new_n3181_ & new_n1941_;
  assign new_n3273_ = ~new_n3215_ | ~new_n3149_;
  assign new_n3274_ = new_n1935_ & new_n3181_ & new_n1941_;
  assign new_n3275_ = ~new_n3216_ | ~new_n3150_;
  assign new_n3276_ = new_n3181_ & new_n1941_;
  assign new_n3277_ = ~new_n3217_ | ~new_n3153_;
  assign new_n3278_ = ~new_n3220_ | ~new_n3156_;
  assign new_n3279_ = ~new_n3221_ | ~new_n3157_;
  assign new_n3280_ = ~new_n2206_ | ~new_n3207_;
  assign new_n3281_ = ~new_n2209_ | ~new_n3209_;
  assign new_n3282_ = new_n2210_ & new_n3210_;
  assign new_n3283_ = new_n1952_ & new_n1955_ & new_n1984_ & new_n3210_ & new_n1962_;
  assign new_n3284_ = ~new_n3222_ | ~new_n3159_;
  assign new_n3285_ = new_n1955_ & new_n1984_ & new_n3210_ & new_n1962_;
  assign new_n3286_ = new_n1955_ & new_n3210_ & new_n1962_;
  assign new_n3287_ = ~new_n3223_ | ~new_n3160_;
  assign new_n3288_ = new_n3210_ & new_n1962_;
  assign new_n3289_ = ~new_n2958_ | ~new_n3238_;
  assign new_n3290_ = ~new_n2960_ | ~new_n3229_;
  assign new_n3291_ = new_n3225_ | new_n3168_;
  assign new_n3292_ = ~new_n2971_ | ~new_n3232_;
  assign new_n3293_ = ~new_n2976_ | ~new_n3227_;
  assign new_n3294_ = ~new_n2843_ | ~new_n3228_;
  assign new_n3295_ = ~new_n2979_ | ~new_n3234_;
  assign new_n3296_ = ~new_n3240_;
  assign new_n3297_ = ~new_n3241_ | ~new_n3176_;
  assign new_n3298_ = ~new_n3242_ | ~new_n3177_;
  assign new_n3299_ = ~new_n3243_ | ~new_n3178_;
  assign new_n3300_ = ~new_n3244_ | ~new_n3180_;
  assign new_n3301_ = ~new_n3245_;
  assign new_n3302_ = ~new_n2670_ | ~new_n3249_;
  assign new_n3303_ = ~new_n2671_ | ~new_n3250_;
  assign new_n3304_ = new_n2374_ & new_n3254_;
  assign new_n3305_ = new_n2082_ & new_n2087_ & new_n2085_ & new_n3254_ & new_n2088_;
  assign new_n3306_ = new_n2087_ & new_n2085_ & new_n3254_ & new_n2088_;
  assign new_n3307_ = ~new_n3251_ | ~new_n3187_;
  assign new_n3308_ = ~new_n3252_ | ~new_n3188_;
  assign new_n3309_ = new_n2087_ & new_n3254_ & new_n2088_;
  assign new_n3310_ = new_n3254_ & new_n2088_;
  assign new_n3311_ = ~new_n3253_;
  assign new_n3312_ = new_n3254_;
  assign new_n3313_ = ~new_n2720_ | ~new_n3258_;
  assign new_n3314_ = ~new_n2721_ | ~new_n3259_;
  assign po065 = new_n3261_ | new_n3199_;
  assign po066 = new_n3262_ | new_n3200_;
  assign new_n3317_ = ~new_n2920_ | ~new_n3296_;
  assign new_n3318_ = ~new_n3264_ | ~new_n3205_;
  assign new_n3319_ = ~new_n3266_;
  assign new_n3320_ = ~new_n3267_;
  assign new_n3321_ = ~new_n3268_ | ~new_n3211_;
  assign new_n3322_ = ~new_n3269_ | ~new_n3212_;
  assign new_n3323_ = new_n2520_ | new_n3270_;
  assign new_n3324_ = ~new_n3273_ | ~new_n2778_;
  assign new_n3325_ = ~new_n3275_ | ~new_n2779_;
  assign new_n3326_ = new_n3271_ | new_n2195_ | new_n2181_ | new_n1004_ | new_n2168_;
  assign new_n3327_ = new_n3272_ | new_n2198_ | new_n1009_ | new_n2183_;
  assign new_n3328_ = ~new_n3273_;
  assign new_n3329_ = new_n3274_ | new_n1014_ | new_n2197_;
  assign new_n3330_ = ~new_n3275_;
  assign new_n3331_ = new_n1019_ | new_n3276_;
  assign new_n3332_ = ~new_n3245_ | ~new_n2539_;
  assign new_n3333_ = ~new_n3279_ | ~new_n1307_;
  assign new_n3334_ = ~new_n3278_ | ~new_n1310_;
  assign new_n3335_ = ~new_n3278_;
  assign new_n3336_ = ~new_n3279_;
  assign new_n3337_ = new_n2792_ & new_n3281_;
  assign new_n3338_ = new_n2543_ | new_n3282_;
  assign new_n3339_ = new_n2793_ & new_n3280_;
  assign new_n3340_ = ~new_n3284_ | ~new_n2794_;
  assign new_n3341_ = ~new_n3287_ | ~new_n2795_;
  assign new_n3342_ = new_n3283_ | new_n2240_ | new_n2224_ | new_n1039_ | new_n2273_;
  assign new_n3343_ = ~new_n3284_;
  assign new_n3344_ = new_n3286_ | new_n1044_ | new_n2242_;
  assign new_n3345_ = ~new_n3287_;
  assign new_n3346_ = new_n1049_ | new_n3288_;
  assign new_n3347_ = ~new_n3267_ | ~new_n2564_;
  assign new_n3348_ = ~new_n3289_ | ~new_n3224_;
  assign new_n3349_ = ~new_n3290_ | ~new_n3226_;
  assign new_n3350_ = ~new_n2584_ | ~new_n3291_;
  assign new_n3351_ = new_n3285_ | new_n2243_ | new_n1090_ | new_n2226_;
  assign new_n3352_ = ~new_n3292_ | ~new_n3233_;
  assign new_n3353_ = ~new_n3293_ | ~new_n3235_;
  assign new_n3354_ = ~new_n3294_ | ~new_n3236_;
  assign new_n3355_ = ~new_n3295_ | ~new_n3237_;
  assign new_n3356_ = ~new_n3302_ | ~new_n3247_;
  assign new_n3357_ = ~new_n3303_ | ~new_n3248_;
  assign new_n3358_ = new_n2687_ | new_n3304_;
  assign new_n3359_ = new_n3305_ | new_n2403_ | new_n2391_ | new_n1228_ | new_n2382_;
  assign new_n3360_ = ~new_n3307_ | ~new_n2883_;
  assign new_n3361_ = ~new_n3308_ | ~new_n2884_;
  assign new_n3362_ = new_n3306_ | new_n2406_ | new_n1230_ | new_n2393_;
  assign new_n3363_ = new_n3309_ | new_n1232_ | new_n2405_;
  assign new_n3364_ = ~new_n3307_;
  assign new_n3365_ = ~new_n3308_;
  assign new_n3366_ = new_n1234_ | new_n3310_;
  assign new_n3367_ = ~new_n3312_ | ~new_n2707_;
  assign new_n3368_ = ~new_n3312_;
  assign new_n3369_ = ~new_n3313_ | ~new_n3255_;
  assign new_n3370_ = ~new_n3314_ | ~new_n3256_;
  assign new_n3371_ = ~new_n3318_ | ~new_n2914_;
  assign new_n3372_ = ~new_n3317_ | ~new_n3263_;
  assign new_n3373_ = ~new_n3318_;
  assign new_n3374_ = new_n3355_ & new_n3352_ & new_n3277_ & new_n3265_;
  assign new_n3375_ = new_n3323_ & new_n3051_;
  assign new_n3376_ = new_n3323_ & new_n3054_;
  assign new_n3377_ = ~new_n3321_;
  assign new_n3378_ = ~new_n3322_;
  assign new_n3379_ = new_n3323_ & new_n2146_;
  assign new_n3380_ = new_n3323_ & new_n3056_;
  assign new_n3381_ = ~new_n3321_ | ~new_n2510_;
  assign new_n3382_ = ~new_n3322_ | ~new_n2511_;
  assign new_n3383_ = ~new_n3323_;
  assign new_n3384_ = ~new_n3326_ | ~new_n2521_;
  assign new_n3385_ = ~new_n2522_ | ~new_n3328_;
  assign new_n3386_ = ~new_n2523_ | ~new_n3330_;
  assign new_n3387_ = ~new_n3326_;
  assign new_n3388_ = ~new_n3327_ | ~new_n2524_;
  assign new_n3389_ = ~new_n3327_;
  assign new_n3390_ = ~new_n3329_ | ~new_n2532_;
  assign new_n3391_ = ~new_n3329_;
  assign new_n3392_ = ~new_n3331_ | ~new_n2534_;
  assign new_n3393_ = ~new_n3331_;
  assign new_n3394_ = ~new_n2203_ | ~new_n3301_;
  assign new_n3395_ = new_n3337_ & new_n1301_;
  assign new_n3396_ = new_n1947_ & new_n3338_;
  assign new_n3397_ = ~new_n1028_ | ~new_n3336_;
  assign new_n3398_ = ~new_n1029_ | ~new_n3335_;
  assign new_n3399_ = new_n3338_ & new_n1314_;
  assign new_n3400_ = ~new_n3337_;
  assign new_n3401_ = ~new_n3338_;
  assign new_n3402_ = ~new_n3339_;
  assign new_n3403_ = ~new_n3342_ | ~new_n2551_;
  assign new_n3404_ = ~new_n2552_ | ~new_n3343_;
  assign new_n3405_ = ~new_n2553_ | ~new_n3345_;
  assign new_n3406_ = ~new_n3342_;
  assign new_n3407_ = ~new_n3351_ | ~new_n2554_;
  assign new_n3408_ = ~new_n3344_;
  assign new_n3409_ = ~new_n3346_ | ~new_n2558_;
  assign new_n3410_ = ~new_n3346_;
  assign new_n3411_ = ~new_n2248_ | ~new_n3320_;
  assign new_n3412_ = ~new_n3351_;
  assign new_n3413_ = ~new_n3344_ | ~new_n2594_;
  assign new_n3414_ = new_n2980_ & new_n3350_;
  assign new_n3415_ = new_n3339_ & new_n1807_;
  assign new_n3416_ = new_n3338_ & new_n2310_;
  assign new_n3417_ = new_n3348_ & new_n3354_ & new_n3297_ & new_n3298_;
  assign new_n3418_ = new_n3349_ & new_n3353_ & new_n3300_ & new_n3299_;
  assign new_n3419_ = new_n2071_ & new_n3402_;
  assign new_n3420_ = new_n3358_ & new_n3106_;
  assign new_n3421_ = ~new_n3356_;
  assign new_n3422_ = ~new_n3357_;
  assign new_n3423_ = new_n3358_ & new_n3110_;
  assign new_n3424_ = ~new_n3356_ | ~new_n2684_;
  assign new_n3425_ = ~new_n3357_ | ~new_n2685_;
  assign new_n3426_ = new_n3358_ & new_n2370_;
  assign new_n3427_ = new_n3358_ & new_n3113_;
  assign new_n3428_ = ~new_n3358_;
  assign new_n3429_ = ~new_n3359_ | ~new_n2692_;
  assign new_n3430_ = ~new_n3359_;
  assign new_n3431_ = ~new_n2693_ | ~new_n3364_;
  assign new_n3432_ = ~new_n2694_ | ~new_n3365_;
  assign new_n3433_ = ~new_n3362_ | ~new_n2695_;
  assign new_n3434_ = ~new_n3362_;
  assign new_n3435_ = ~new_n3363_ | ~new_n2702_;
  assign new_n3436_ = ~new_n3363_;
  assign new_n3437_ = ~new_n3366_ | ~new_n2706_;
  assign new_n3438_ = ~new_n3366_;
  assign new_n3439_ = ~new_n2413_ | ~new_n3368_;
  assign new_n3440_ = ~new_n3369_;
  assign new_n3441_ = ~new_n3370_;
  assign new_n3442_ = ~new_n3369_ | ~new_n2734_;
  assign new_n3443_ = ~new_n3370_ | ~new_n2735_;
  assign new_n3444_ = ~new_n2744_ | ~new_n3373_;
  assign new_n3445_ = ~new_n3372_ | ~new_n3042_;
  assign new_n3446_ = ~new_n3372_;
  assign po070 = ~new_n3374_;
  assign new_n3448_ = new_n3417_ & new_n3418_ & new_n3374_;
  assign new_n3449_ = new_n3140_ & new_n3383_;
  assign new_n3450_ = new_n3145_ & new_n3383_;
  assign new_n3451_ = new_n2933_ & new_n3383_;
  assign new_n3452_ = new_n1921_ & new_n3383_;
  assign new_n3453_ = ~new_n2147_ | ~new_n3377_;
  assign new_n3454_ = ~new_n2148_ | ~new_n3378_;
  assign new_n3455_ = ~new_n2157_ | ~new_n3387_;
  assign new_n3456_ = ~new_n3385_ | ~new_n3324_;
  assign new_n3457_ = ~new_n3386_ | ~new_n3325_;
  assign new_n3458_ = ~new_n2160_ | ~new_n3389_;
  assign new_n3459_ = ~new_n2175_ | ~new_n3391_;
  assign new_n3460_ = ~new_n2184_ | ~new_n3393_;
  assign po073 = ~new_n3394_ | ~new_n3332_;
  assign new_n3462_ = new_n1945_ & new_n3400_;
  assign new_n3463_ = new_n1302_ & new_n3401_;
  assign new_n3464_ = ~new_n3397_ | ~new_n3333_;
  assign new_n3465_ = ~new_n3398_ | ~new_n3334_;
  assign new_n3466_ = new_n1032_ & new_n3401_;
  assign new_n3467_ = ~new_n2211_ | ~new_n3406_;
  assign new_n3468_ = ~new_n3404_ | ~new_n3340_;
  assign new_n3469_ = ~new_n3405_ | ~new_n3341_;
  assign new_n3470_ = ~new_n2214_ | ~new_n3412_;
  assign new_n3471_ = ~new_n2227_ | ~new_n3410_;
  assign po074 = ~new_n3411_ | ~new_n3347_;
  assign new_n3473_ = ~new_n2277_ | ~new_n3408_;
  assign new_n3474_ = new_n3414_ & new_n2842_;
  assign new_n3475_ = ~new_n3414_;
  assign new_n3476_ = new_n2036_ & new_n3401_;
  assign po071 = ~new_n3417_;
  assign po069 = ~new_n3418_;
  assign new_n3479_ = new_n3183_ & new_n3428_;
  assign new_n3480_ = new_n3184_ & new_n3428_;
  assign new_n3481_ = new_n3015_ & new_n3428_;
  assign new_n3482_ = ~new_n2368_ | ~new_n3421_;
  assign new_n3483_ = ~new_n2369_ | ~new_n3422_;
  assign new_n3484_ = new_n2079_ & new_n3428_;
  assign new_n3485_ = ~new_n2375_ | ~new_n3430_;
  assign new_n3486_ = ~new_n3431_ | ~new_n3360_;
  assign new_n3487_ = ~new_n3432_ | ~new_n3361_;
  assign new_n3488_ = ~new_n2378_ | ~new_n3434_;
  assign new_n3489_ = ~new_n2390_ | ~new_n3436_;
  assign new_n3490_ = ~new_n2402_ | ~new_n3438_;
  assign po091 = ~new_n3439_ | ~new_n3367_;
  assign new_n3492_ = ~new_n2451_ | ~new_n3440_;
  assign new_n3493_ = ~new_n2452_ | ~new_n3441_;
  assign new_n3494_ = ~new_n3444_ | ~new_n3371_;
  assign new_n3495_ = ~new_n2915_ | ~new_n3446_;
  assign po087 = new_n3449_ | new_n3375_;
  assign po088 = new_n3450_ | new_n3376_;
  assign po090 = new_n3452_ | new_n3379_;
  assign po089 = new_n3451_ | new_n3380_;
  assign new_n3500_ = ~new_n3453_ | ~new_n3381_;
  assign new_n3501_ = ~new_n3454_ | ~new_n3382_;
  assign po077 = ~new_n3455_ | ~new_n3384_;
  assign new_n3503_ = ~new_n3456_;
  assign new_n3504_ = ~new_n3457_;
  assign po078 = ~new_n3458_ | ~new_n3388_;
  assign po079 = ~new_n3459_ | ~new_n3390_;
  assign po080 = ~new_n3460_ | ~new_n3392_;
  assign new_n3508_ = ~new_n3456_ | ~new_n2537_;
  assign new_n3509_ = ~new_n3457_ | ~new_n2538_;
  assign po076 = new_n3462_ | new_n3395_;
  assign po086 = new_n3463_ | new_n3396_;
  assign new_n3512_ = new_n3466_ | new_n3399_;
  assign new_n3513_ = new_n3319_ & new_n3464_ & new_n2542_;
  assign new_n3514_ = new_n3319_ & new_n3465_ & new_n2792_;
  assign new_n3515_ = new_n3266_ & new_n3465_ & new_n2948_;
  assign new_n3516_ = new_n3266_ & new_n3464_ & new_n3067_;
  assign po081 = ~new_n3467_ | ~new_n3403_;
  assign new_n3518_ = ~new_n3468_;
  assign new_n3519_ = ~new_n3469_;
  assign po082 = ~new_n3470_ | ~new_n3407_;
  assign po084 = ~new_n3471_ | ~new_n3409_;
  assign new_n3522_ = ~new_n3468_ | ~new_n2562_;
  assign new_n3523_ = ~new_n3469_ | ~new_n2563_;
  assign new_n3524_ = new_n3448_ & new_n498_ & new_n495_;
  assign po083 = ~new_n3473_ | ~new_n3413_;
  assign new_n3526_ = new_n3083_ & new_n3475_;
  assign po072 = new_n3419_ | new_n3415_;
  assign new_n3528_ = new_n3476_ | new_n3416_;
  assign po100 = new_n3479_ | new_n3420_;
  assign po101 = new_n3480_ | new_n3423_;
  assign new_n3531_ = ~new_n3482_ | ~new_n3424_;
  assign new_n3532_ = ~new_n3483_ | ~new_n3425_;
  assign po103 = new_n3484_ | new_n3426_;
  assign po102 = new_n3481_ | new_n3427_;
  assign po096 = ~new_n3485_ | ~new_n3429_;
  assign new_n3536_ = ~new_n3486_;
  assign new_n3537_ = ~new_n3487_;
  assign po097 = ~new_n3488_ | ~new_n3433_;
  assign po098 = ~new_n3489_ | ~new_n3435_;
  assign po099 = ~new_n3490_ | ~new_n3437_;
  assign new_n3541_ = ~new_n3486_ | ~new_n2708_;
  assign new_n3542_ = ~new_n3487_ | ~new_n2709_;
  assign new_n3543_ = ~new_n3492_ | ~new_n3442_;
  assign new_n3544_ = ~new_n3493_ | ~new_n3443_;
  assign new_n3545_ = ~new_n3494_;
  assign new_n3546_ = ~new_n3495_ | ~new_n3445_;
  assign new_n3547_ = ~new_n3501_ | ~new_n2504_;
  assign new_n3548_ = ~new_n3500_ | ~new_n2505_;
  assign new_n3549_ = ~new_n3500_;
  assign new_n3550_ = ~new_n3501_;
  assign new_n3551_ = ~new_n2199_ | ~new_n3503_;
  assign new_n3552_ = ~new_n2200_ | ~new_n3504_;
  assign po094 = new_n3512_;
  assign po095 = new_n3512_;
  assign new_n3555_ = new_n3516_ | new_n3515_ | new_n3514_ | new_n3513_;
  assign new_n3556_ = ~new_n2244_ | ~new_n3518_;
  assign new_n3557_ = ~new_n2245_ | ~new_n3519_;
  assign po085 = ~new_n3524_;
  assign po075 = new_n3526_ | new_n3474_;
  assign po092 = new_n3528_;
  assign po093 = new_n3528_;
  assign new_n3562_ = ~new_n3494_ | ~new_n2989_;
  assign new_n3563_ = ~new_n3532_ | ~new_n2681_;
  assign new_n3564_ = ~new_n3531_ | ~new_n2682_;
  assign new_n3565_ = ~new_n3531_;
  assign new_n3566_ = ~new_n3532_;
  assign new_n3567_ = ~new_n2414_ | ~new_n3536_;
  assign new_n3568_ = ~new_n2415_ | ~new_n3537_;
  assign new_n3569_ = ~new_n3544_ | ~new_n2729_;
  assign new_n3570_ = ~new_n3543_ | ~new_n2730_;
  assign new_n3571_ = ~new_n3543_;
  assign new_n3572_ = ~new_n3544_;
  assign new_n3573_ = ~new_n3546_;
  assign new_n3574_ = ~new_n2132_ | ~new_n3550_;
  assign new_n3575_ = ~new_n2133_ | ~new_n3549_;
  assign new_n3576_ = ~new_n3551_ | ~new_n3508_;
  assign new_n3577_ = ~new_n3552_ | ~new_n3509_;
  assign new_n3578_ = ~new_n3555_;
  assign new_n3579_ = ~new_n3556_ | ~new_n3522_;
  assign new_n3580_ = ~new_n3557_ | ~new_n3523_;
  assign new_n3581_ = ~new_n2855_ | ~new_n3545_;
  assign new_n3582_ = ~new_n3546_ | ~new_n2990_;
  assign new_n3583_ = ~new_n2357_ | ~new_n3566_;
  assign new_n3584_ = ~new_n2358_ | ~new_n3565_;
  assign new_n3585_ = ~new_n3567_ | ~new_n3541_;
  assign new_n3586_ = ~new_n3568_ | ~new_n3542_;
  assign new_n3587_ = ~new_n2437_ | ~new_n3572_;
  assign new_n3588_ = ~new_n2438_ | ~new_n3571_;
  assign new_n3589_ = ~new_n3574_ | ~new_n3547_;
  assign new_n3590_ = ~new_n3575_ | ~new_n3548_;
  assign new_n3591_ = ~new_n3577_ | ~new_n2535_;
  assign new_n3592_ = ~new_n3576_ | ~new_n2536_;
  assign new_n3593_ = ~new_n3576_;
  assign new_n3594_ = ~new_n3577_;
  assign new_n3595_ = ~new_n3580_ | ~new_n2560_;
  assign new_n3596_ = ~new_n3579_ | ~new_n2561_;
  assign new_n3597_ = ~new_n3579_;
  assign new_n3598_ = ~new_n3580_;
  assign new_n3599_ = ~new_n3581_ | ~new_n3562_;
  assign new_n3600_ = ~new_n2856_ | ~new_n3573_;
  assign new_n3601_ = ~new_n3583_ | ~new_n3563_;
  assign new_n3602_ = ~new_n3584_ | ~new_n3564_;
  assign new_n3603_ = ~new_n3586_ | ~new_n2704_;
  assign new_n3604_ = ~new_n3585_ | ~new_n2705_;
  assign new_n3605_ = ~new_n3585_;
  assign new_n3606_ = ~new_n3586_;
  assign new_n3607_ = ~new_n3587_ | ~new_n3569_;
  assign new_n3608_ = ~new_n3588_ | ~new_n3570_;
  assign new_n3609_ = ~new_n3599_ | ~new_n2756_;
  assign new_n3610_ = ~new_n3590_ | ~new_n2485_;
  assign new_n3611_ = ~new_n3589_ | ~new_n2486_;
  assign new_n3612_ = ~new_n3589_;
  assign new_n3613_ = ~new_n3590_;
  assign new_n3614_ = ~new_n2185_ | ~new_n3594_;
  assign new_n3615_ = ~new_n2186_ | ~new_n3593_;
  assign new_n3616_ = ~new_n2230_ | ~new_n3598_;
  assign new_n3617_ = ~new_n2232_ | ~new_n3597_;
  assign new_n3618_ = ~new_n3599_;
  assign new_n3619_ = ~new_n3600_ | ~new_n3582_;
  assign new_n3620_ = ~new_n3602_ | ~new_n2663_;
  assign new_n3621_ = ~new_n3601_ | ~new_n2664_;
  assign new_n3622_ = ~new_n3601_;
  assign new_n3623_ = ~new_n3602_;
  assign new_n3624_ = ~new_n2399_ | ~new_n3606_;
  assign new_n3625_ = ~new_n2400_ | ~new_n3605_;
  assign new_n3626_ = ~new_n3608_ | ~new_n2713_;
  assign new_n3627_ = ~new_n3607_ | ~new_n2714_;
  assign new_n3628_ = ~new_n3607_;
  assign new_n3629_ = ~new_n3608_;
  assign new_n3630_ = ~new_n3619_ | ~new_n2755_;
  assign new_n3631_ = ~new_n2479_ | ~new_n3618_;
  assign new_n3632_ = ~new_n2109_ | ~new_n3613_;
  assign new_n3633_ = ~new_n2110_ | ~new_n3612_;
  assign new_n3634_ = ~new_n3614_ | ~new_n3591_;
  assign new_n3635_ = ~new_n3615_ | ~new_n3592_;
  assign new_n3636_ = ~new_n3616_ | ~new_n3595_;
  assign new_n3637_ = ~new_n3617_ | ~new_n3596_;
  assign new_n3638_ = ~new_n3619_;
  assign new_n3639_ = ~new_n2334_ | ~new_n3623_;
  assign new_n3640_ = ~new_n2335_ | ~new_n3622_;
  assign new_n3641_ = ~new_n3624_ | ~new_n3603_;
  assign new_n3642_ = ~new_n3625_ | ~new_n3604_;
  assign new_n3643_ = ~new_n2417_ | ~new_n3629_;
  assign new_n3644_ = ~new_n2418_ | ~new_n3628_;
  assign new_n3645_ = ~new_n2478_ | ~new_n3638_;
  assign new_n3646_ = ~new_n3631_ | ~new_n3609_;
  assign new_n3647_ = ~new_n3632_ | ~new_n3610_;
  assign new_n3648_ = ~new_n3633_ | ~new_n3611_;
  assign new_n3649_ = ~new_n3635_ | ~new_n2517_;
  assign new_n3650_ = ~new_n3634_ | ~new_n2518_;
  assign new_n3651_ = ~new_n3634_;
  assign new_n3652_ = ~new_n3635_;
  assign new_n3653_ = ~new_n3637_ | ~new_n2548_;
  assign new_n3654_ = ~new_n3636_ | ~new_n2549_;
  assign new_n3655_ = ~new_n3636_;
  assign new_n3656_ = ~new_n3637_;
  assign new_n3657_ = ~new_n3639_ | ~new_n3620_;
  assign new_n3658_ = ~new_n3640_ | ~new_n3621_;
  assign new_n3659_ = ~new_n3642_ | ~new_n2689_;
  assign new_n3660_ = ~new_n3641_ | ~new_n2690_;
  assign new_n3661_ = ~new_n3641_;
  assign new_n3662_ = ~new_n3642_;
  assign new_n3663_ = ~new_n3643_ | ~new_n3626_;
  assign new_n3664_ = ~new_n3644_ | ~new_n3627_;
  assign new_n3665_ = ~new_n3646_ | ~new_n2741_;
  assign new_n3666_ = ~new_n3645_ | ~new_n3630_;
  assign new_n3667_ = ~new_n3646_;
  assign new_n3668_ = ~new_n3647_;
  assign new_n3669_ = ~new_n3648_;
  assign new_n3670_ = ~new_n3648_ | ~new_n2498_;
  assign new_n3671_ = ~new_n3647_ | ~new_n2499_;
  assign new_n3672_ = ~new_n2153_ | ~new_n3652_;
  assign new_n3673_ = ~new_n2154_ | ~new_n3651_;
  assign new_n3674_ = ~new_n2207_ | ~new_n3656_;
  assign new_n3675_ = ~new_n2208_ | ~new_n3655_;
  assign new_n3676_ = ~new_n3657_;
  assign new_n3677_ = ~new_n3658_;
  assign new_n3678_ = ~new_n3658_ | ~new_n2674_;
  assign new_n3679_ = ~new_n3657_ | ~new_n2675_;
  assign new_n3680_ = ~new_n2371_ | ~new_n3662_;
  assign new_n3681_ = ~new_n2372_ | ~new_n3661_;
  assign new_n3682_ = ~new_n3663_;
  assign new_n3683_ = ~new_n3664_;
  assign new_n3684_ = ~new_n3664_ | ~new_n2724_;
  assign new_n3685_ = ~new_n3663_ | ~new_n2725_;
  assign new_n3686_ = ~new_n2455_ | ~new_n3667_;
  assign new_n3687_ = ~new_n3666_ | ~new_n2742_;
  assign new_n3688_ = ~new_n3666_;
  assign new_n3689_ = ~new_n2120_ | ~new_n3669_;
  assign new_n3690_ = ~new_n2122_ | ~new_n3668_;
  assign new_n3691_ = ~new_n3672_ | ~new_n3649_;
  assign new_n3692_ = ~new_n3673_ | ~new_n3650_;
  assign new_n3693_ = ~new_n3674_ | ~new_n3653_;
  assign new_n3694_ = ~new_n3675_ | ~new_n3654_;
  assign new_n3695_ = ~new_n2344_ | ~new_n3677_;
  assign new_n3696_ = ~new_n2346_ | ~new_n3676_;
  assign new_n3697_ = ~new_n3680_ | ~new_n3659_;
  assign new_n3698_ = ~new_n3681_ | ~new_n3660_;
  assign new_n3699_ = ~new_n2427_ | ~new_n3683_;
  assign new_n3700_ = ~new_n2429_ | ~new_n3682_;
  assign new_n3701_ = ~new_n3686_ | ~new_n3665_;
  assign new_n3702_ = ~new_n2456_ | ~new_n3688_;
  assign new_n3703_ = ~new_n3689_ | ~new_n3670_;
  assign new_n3704_ = ~new_n3690_ | ~new_n3671_;
  assign new_n3705_ = ~new_n3691_;
  assign new_n3706_ = ~new_n3692_;
  assign new_n3707_ = ~new_n3691_ | ~new_n2530_;
  assign new_n3708_ = ~new_n3692_ | ~new_n2531_;
  assign new_n3709_ = ~new_n3693_;
  assign new_n3710_ = ~new_n3694_;
  assign new_n3711_ = ~new_n3693_ | ~new_n2592_;
  assign new_n3712_ = ~new_n3694_ | ~new_n2593_;
  assign new_n3713_ = ~new_n3695_ | ~new_n3678_;
  assign new_n3714_ = ~new_n3696_ | ~new_n3679_;
  assign new_n3715_ = ~new_n3697_;
  assign new_n3716_ = ~new_n3698_;
  assign new_n3717_ = ~new_n3697_ | ~new_n2700_;
  assign new_n3718_ = ~new_n3698_ | ~new_n2701_;
  assign new_n3719_ = ~new_n3699_ | ~new_n3684_;
  assign new_n3720_ = ~new_n3700_ | ~new_n3685_;
  assign new_n3721_ = ~new_n3701_;
  assign new_n3722_ = ~new_n3702_ | ~new_n3687_;
  assign new_n3723_ = ~new_n3701_ | ~new_n2751_;
  assign new_n3724_ = new_n3246_ & new_n3703_ & new_n2516_;
  assign new_n3725_ = new_n3246_ & new_n3704_ & new_n2777_;
  assign new_n3726_ = new_n3182_ & new_n3704_ & new_n2937_;
  assign new_n3727_ = new_n3182_ & new_n3703_ & new_n3059_;
  assign new_n3728_ = ~new_n2172_ | ~new_n3705_;
  assign new_n3729_ = ~new_n2173_ | ~new_n3706_;
  assign new_n3730_ = ~new_n2275_ | ~new_n3709_;
  assign new_n3731_ = ~new_n2276_ | ~new_n3710_;
  assign new_n3732_ = new_n317_ & new_n3720_ & new_n3039_;
  assign new_n3733_ = new_n317_ & new_n3719_ & new_n3128_;
  assign new_n3734_ = new_n426_ & new_n3720_ & new_n2911_;
  assign new_n3735_ = new_n426_ & new_n3719_ & new_n2738_;
  assign new_n3736_ = new_n3311_ & new_n3713_ & new_n2688_;
  assign new_n3737_ = new_n3311_ & new_n3714_ & new_n2882_;
  assign new_n3738_ = new_n3253_ & new_n3714_ & new_n3019_;
  assign new_n3739_ = new_n3253_ & new_n3713_ & new_n3114_;
  assign new_n3740_ = ~new_n2387_ | ~new_n3715_;
  assign new_n3741_ = ~new_n2388_ | ~new_n3716_;
  assign new_n3742_ = ~new_n3722_;
  assign new_n3743_ = ~new_n2468_ | ~new_n3721_;
  assign new_n3744_ = ~new_n3722_ | ~new_n2752_;
  assign new_n3745_ = new_n3727_ | new_n3726_ | new_n3725_ | new_n3724_;
  assign new_n3746_ = ~new_n3728_ | ~new_n3707_;
  assign new_n3747_ = ~new_n3729_ | ~new_n3708_;
  assign new_n3748_ = ~new_n3730_ | ~new_n3711_;
  assign new_n3749_ = ~new_n3731_ | ~new_n3712_;
  assign new_n3750_ = new_n3733_ | new_n3732_ | new_n3734_ | new_n3735_;
  assign new_n3751_ = new_n3739_ | new_n3738_ | new_n3737_ | new_n3736_;
  assign new_n3752_ = ~new_n3740_ | ~new_n3717_;
  assign new_n3753_ = ~new_n3741_ | ~new_n3718_;
  assign new_n3754_ = ~new_n3743_ | ~new_n3723_;
  assign new_n3755_ = ~new_n2469_ | ~new_n3742_;
  assign new_n3756_ = ~new_n3745_;
  assign new_n3757_ = ~new_n3746_ | ~new_n2525_;
  assign new_n3758_ = ~new_n3747_ | ~new_n2526_;
  assign new_n3759_ = ~new_n3746_;
  assign new_n3760_ = ~new_n3747_;
  assign new_n3761_ = ~new_n3748_ | ~new_n2555_;
  assign new_n3762_ = ~new_n3749_ | ~new_n2556_;
  assign new_n3763_ = ~new_n3748_;
  assign new_n3764_ = ~new_n3749_;
  assign new_n3765_ = ~new_n3750_;
  assign new_n3766_ = ~new_n3751_;
  assign new_n3767_ = ~new_n3752_ | ~new_n2696_;
  assign new_n3768_ = ~new_n3753_ | ~new_n2697_;
  assign new_n3769_ = ~new_n3752_;
  assign new_n3770_ = ~new_n3753_;
  assign new_n3771_ = ~new_n3754_ | ~new_n2745_;
  assign new_n3772_ = ~new_n3754_;
  assign new_n3773_ = ~new_n3755_ | ~new_n3744_;
  assign new_n3774_ = ~new_n2161_ | ~new_n3759_;
  assign new_n3775_ = ~new_n2163_ | ~new_n3760_;
  assign new_n3776_ = ~new_n2215_ | ~new_n3763_;
  assign new_n3777_ = ~new_n2217_ | ~new_n3764_;
  assign new_n3778_ = ~new_n2379_ | ~new_n3769_;
  assign new_n3779_ = ~new_n2381_ | ~new_n3770_;
  assign new_n3780_ = ~new_n2459_ | ~new_n3772_;
  assign new_n3781_ = ~new_n3773_ | ~new_n2747_;
  assign new_n3782_ = ~new_n3773_;
  assign new_n3783_ = ~new_n3774_ | ~new_n3757_;
  assign new_n3784_ = ~new_n3775_ | ~new_n3758_;
  assign new_n3785_ = ~new_n3776_ | ~new_n3761_;
  assign new_n3786_ = ~new_n3777_ | ~new_n3762_;
  assign new_n3787_ = new_n3182_ & new_n3784_;
  assign new_n3788_ = ~new_n3778_ | ~new_n3767_;
  assign new_n3789_ = ~new_n3779_ | ~new_n3768_;
  assign new_n3790_ = ~new_n3780_ | ~new_n3771_;
  assign new_n3791_ = ~new_n2460_ | ~new_n3782_;
  assign new_n3792_ = new_n3266_ & new_n3786_;
  assign new_n3793_ = ~new_n3783_;
  assign new_n3794_ = ~new_n3785_;
  assign new_n3795_ = new_n3793_ & new_n3246_;
  assign new_n3796_ = ~new_n3788_;
  assign new_n3797_ = new_n3253_ & new_n3789_;
  assign new_n3798_ = ~new_n3790_;
  assign new_n3799_ = ~new_n3791_ | ~new_n3781_;
  assign new_n3800_ = new_n3794_ & new_n3319_;
  assign new_n3801_ = new_n317_ & new_n3799_;
  assign new_n3802_ = new_n3798_ & new_n426_;
  assign new_n3803_ = new_n3795_ | new_n3787_;
  assign new_n3804_ = new_n3796_ & new_n3311_;
  assign new_n3805_ = new_n3800_ | new_n3792_;
  assign new_n3806_ = new_n3802_ | new_n3801_;
  assign new_n3807_ = ~new_n3803_;
  assign new_n3808_ = new_n3804_ | new_n3797_;
  assign new_n3809_ = ~new_n3805_;
  assign new_n3810_ = ~new_n3803_ | ~new_n3756_;
  assign new_n3811_ = ~new_n3805_ | ~new_n3578_;
  assign new_n3812_ = ~new_n3806_ | ~new_n3765_;
  assign new_n3813_ = ~new_n3806_;
  assign new_n3814_ = ~new_n3808_ | ~new_n3766_;
  assign new_n3815_ = ~new_n3808_;
  assign new_n3816_ = ~new_n3745_ | ~new_n3807_;
  assign new_n3817_ = ~new_n3555_ | ~new_n3809_;
  assign new_n3818_ = ~new_n3750_ | ~new_n3813_;
  assign new_n3819_ = ~new_n3751_ | ~new_n3815_;
  assign new_n3820_ = ~new_n3810_ | ~new_n3816_;
  assign new_n3821_ = ~new_n3811_ | ~new_n3817_;
  assign new_n3822_ = ~new_n3812_ | ~new_n3818_;
  assign new_n3823_ = ~new_n3814_ | ~new_n3819_;
  assign po104 = ~new_n3820_;
  assign po105 = ~new_n3821_;
  assign po107 = ~new_n3822_;
  assign po106 = ~new_n3823_;
  assign po000 = pi164;
endmodule


