// Benchmark "i3" written by ABC on Thu Mar 19 13:02:36 2020

module i3 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131,
    po0, po1, po2, po3, po4, po5  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131;
  output po0, po1, po2, po3, po4, po5;
  wire new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_,
    new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_,
    new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_,
    new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_,
    new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n203_, new_n204_;
  assign po0 = pi000 | pi001;
  assign po1 = pi002 | pi003;
  assign new_n141_ = pi004 | pi005;
  assign new_n142_ = pi006 | pi007;
  assign new_n143_ = pi008 | pi009;
  assign new_n144_ = pi010 | pi011;
  assign new_n145_ = pi012 | pi013;
  assign new_n146_ = pi014 | pi015;
  assign new_n147_ = pi016 | pi017;
  assign new_n148_ = pi018 | pi019;
  assign new_n149_ = pi020 | pi021;
  assign new_n150_ = pi022 | pi023;
  assign new_n151_ = pi024 | pi025;
  assign new_n152_ = pi026 | pi027;
  assign new_n153_ = pi028 | pi029;
  assign new_n154_ = pi030 | pi031;
  assign new_n155_ = pi032 | pi033;
  assign new_n156_ = pi034 | pi035;
  assign new_n157_ = pi036 | pi037;
  assign new_n158_ = pi038 | pi039;
  assign new_n159_ = pi040 | pi041;
  assign new_n160_ = pi042 | pi043;
  assign new_n161_ = pi044 | pi045;
  assign new_n162_ = pi046 | pi047;
  assign new_n163_ = pi048 | pi049;
  assign new_n164_ = pi050 | pi051;
  assign new_n165_ = pi052 | pi053;
  assign new_n166_ = pi054 | pi055;
  assign new_n167_ = pi056 | pi057;
  assign new_n168_ = pi058 | pi059;
  assign new_n169_ = pi060 | pi061;
  assign new_n170_ = pi062 | pi063;
  assign new_n171_ = pi064 | pi065;
  assign new_n172_ = pi066 | pi067;
  assign new_n173_ = pi068 | pi069;
  assign new_n174_ = pi070 | pi071;
  assign new_n175_ = pi072 | pi073;
  assign new_n176_ = pi074 | pi075;
  assign new_n177_ = pi076 | pi077;
  assign new_n178_ = pi078 | pi079;
  assign new_n179_ = pi080 | pi081;
  assign new_n180_ = pi082 | pi083;
  assign new_n181_ = pi084 | pi085;
  assign new_n182_ = pi086 | pi087;
  assign new_n183_ = pi088 | pi089;
  assign new_n184_ = pi090 | pi091;
  assign new_n185_ = pi092 | pi093;
  assign new_n186_ = pi094 | pi095;
  assign new_n187_ = pi096 | pi097;
  assign new_n188_ = pi098 | pi099;
  assign new_n189_ = pi100 | pi101;
  assign new_n190_ = pi102 | pi103;
  assign new_n191_ = pi104 | pi105;
  assign new_n192_ = pi106 | pi107;
  assign new_n193_ = pi108 | pi109;
  assign new_n194_ = pi110 | pi111;
  assign new_n195_ = pi112 | pi113;
  assign new_n196_ = pi114 | pi115;
  assign new_n197_ = pi116 | pi117;
  assign new_n198_ = pi118 | pi119;
  assign new_n199_ = pi120 | pi121;
  assign new_n200_ = pi122 | pi123;
  assign new_n201_ = pi124 | pi125;
  assign new_n202_ = pi126 | pi127;
  assign new_n203_ = pi128 | pi129;
  assign new_n204_ = pi130 | pi131;
  assign po2 = new_n152_ & new_n151_ & new_n149_ & new_n150_ & new_n148_ & new_n146_ & new_n145_ & new_n147_ & new_n142_ & new_n141_ & new_n143_ & new_n144_ & new_n154_ & new_n153_ & new_n156_ & new_n155_;
  assign po3 = new_n168_ & new_n167_ & new_n165_ & new_n166_ & new_n164_ & new_n162_ & new_n161_ & new_n163_ & new_n158_ & new_n157_ & new_n159_ & new_n160_ & new_n170_ & new_n169_ & new_n172_ & new_n171_;
  assign po4 = new_n184_ & new_n183_ & new_n181_ & new_n182_ & new_n180_ & new_n178_ & new_n177_ & new_n179_ & new_n174_ & new_n173_ & new_n175_ & new_n176_ & new_n186_ & new_n185_ & new_n188_ & new_n187_;
  assign po5 = new_n200_ & new_n199_ & new_n197_ & new_n198_ & new_n196_ & new_n194_ & new_n193_ & new_n195_ & new_n190_ & new_n189_ & new_n191_ & new_n192_ & new_n202_ & new_n201_ & new_n204_ & new_n203_;
endmodule


