// Benchmark "DES" written by ABC on Thu Mar 19 13:02:36 2020

module DES ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244;
  wire new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_,
    new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_,
    new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_,
    new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_,
    new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_,
    new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_,
    new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_,
    new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_,
    new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_,
    new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_,
    new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_,
    new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_,
    new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_,
    new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_,
    new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_,
    new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_,
    new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_,
    new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_,
    new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_,
    new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_,
    new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_,
    new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_,
    new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_,
    new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_,
    new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_,
    new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_,
    new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_,
    new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_,
    new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_,
    new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_,
    new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_,
    new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_,
    new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_,
    new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_,
    new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_,
    new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_,
    new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_,
    new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_,
    new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_,
    new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_,
    new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_,
    new_n1425_, new_n1426_, new_n1427_;
  assign po000 = new_n1192_;
  assign po001 = new_n1193_;
  assign po002 = new_n1194_;
  assign po003 = new_n1195_;
  assign po004 = new_n1196_;
  assign po005 = new_n1197_;
  assign po006 = new_n1198_;
  assign po007 = new_n1199_;
  assign po008 = new_n1200_;
  assign po009 = new_n1201_;
  assign po010 = new_n1202_;
  assign po011 = new_n1203_;
  assign po012 = new_n1204_;
  assign po013 = new_n1205_;
  assign po014 = new_n1206_;
  assign po015 = new_n1207_;
  assign po016 = new_n1208_;
  assign po017 = new_n1209_;
  assign po018 = new_n1210_;
  assign po019 = new_n1211_;
  assign po020 = new_n1212_;
  assign po021 = new_n1213_;
  assign po022 = new_n1214_;
  assign po023 = new_n1215_;
  assign po024 = new_n1216_;
  assign po025 = new_n1217_;
  assign po026 = new_n1218_;
  assign po027 = new_n1219_;
  assign po028 = new_n1220_;
  assign po029 = new_n1221_;
  assign po030 = new_n1222_;
  assign po031 = new_n1223_;
  assign po032 = new_n1224_;
  assign po033 = new_n1225_;
  assign po034 = new_n1226_;
  assign po035 = new_n1227_;
  assign po036 = new_n1228_;
  assign po037 = new_n1229_;
  assign po038 = new_n1230_;
  assign po039 = new_n1231_;
  assign po040 = new_n1232_;
  assign po041 = new_n1233_;
  assign po042 = new_n1234_;
  assign po043 = new_n1235_;
  assign po044 = new_n1236_;
  assign po045 = new_n1237_;
  assign po046 = new_n1238_;
  assign po047 = new_n1239_;
  assign po048 = new_n1240_;
  assign po049 = new_n1241_;
  assign po050 = new_n1242_;
  assign po051 = new_n1243_;
  assign po052 = new_n1244_;
  assign po053 = new_n1245_;
  assign po054 = new_n1246_;
  assign po055 = new_n1247_;
  assign po056 = new_n750_;
  assign po057 = new_n1322_;
  assign po058 = new_n751_;
  assign po059 = new_n1316_;
  assign po060 = new_n752_;
  assign po061 = new_n1310_;
  assign po062 = new_n753_;
  assign po063 = new_n1285_;
  assign po064 = new_n754_;
  assign po065 = new_n1359_;
  assign po066 = new_n755_;
  assign po067 = new_n1294_;
  assign po068 = new_n756_;
  assign po069 = new_n1355_;
  assign po070 = new_n757_;
  assign po071 = new_n1353_;
  assign po072 = new_n758_;
  assign po073 = new_n1352_;
  assign po074 = new_n759_;
  assign po075 = new_n1351_;
  assign po076 = new_n760_;
  assign po077 = new_n1349_;
  assign po078 = new_n761_;
  assign po079 = new_n1347_;
  assign po080 = new_n762_;
  assign po081 = new_n1345_;
  assign po082 = new_n763_;
  assign po083 = new_n1343_;
  assign po084 = new_n764_;
  assign po085 = new_n1341_;
  assign po086 = new_n765_;
  assign po087 = new_n1339_;
  assign po088 = new_n766_;
  assign po089 = new_n1337_;
  assign po090 = new_n767_;
  assign po091 = new_n1335_;
  assign po092 = new_n768_;
  assign po093 = new_n1333_;
  assign po094 = new_n769_;
  assign po095 = new_n1331_;
  assign po096 = new_n770_;
  assign po097 = new_n1329_;
  assign po098 = new_n771_;
  assign po099 = new_n1327_;
  assign po100 = new_n772_;
  assign po101 = new_n1325_;
  assign po102 = new_n773_;
  assign po103 = new_n1323_;
  assign po104 = new_n774_;
  assign po105 = new_n1321_;
  assign po106 = new_n775_;
  assign po107 = new_n1319_;
  assign po108 = new_n776_;
  assign po109 = new_n1317_;
  assign po110 = new_n777_;
  assign po111 = new_n1315_;
  assign po112 = new_n778_;
  assign po113 = new_n1313_;
  assign po114 = new_n779_;
  assign po115 = new_n1311_;
  assign po116 = new_n780_;
  assign po117 = new_n1309_;
  assign po118 = new_n781_;
  assign po119 = new_n1307_;
  assign po120 = new_n782_;
  assign po121 = new_n783_;
  assign po122 = new_n784_;
  assign po123 = new_n785_;
  assign po124 = new_n786_;
  assign po125 = new_n787_;
  assign po126 = new_n788_;
  assign po127 = new_n789_;
  assign po128 = new_n790_;
  assign po129 = new_n791_;
  assign po130 = new_n792_;
  assign po131 = new_n793_;
  assign po132 = new_n794_;
  assign po133 = new_n810_;
  assign po134 = new_n809_;
  assign po135 = new_n808_;
  assign po136 = new_n807_;
  assign po137 = new_n806_;
  assign po138 = new_n805_;
  assign po139 = new_n804_;
  assign po140 = new_n803_;
  assign po141 = new_n802_;
  assign po142 = new_n801_;
  assign po143 = new_n747_;
  assign po144 = new_n748_;
  assign po145 = new_n749_;
  assign po146 = new_n795_;
  assign po147 = new_n796_;
  assign po148 = new_n797_;
  assign po149 = new_n798_;
  assign po150 = new_n799_;
  assign po151 = new_n800_;
  assign po152 = new_n1279_;
  assign po153 = new_n1278_;
  assign po154 = new_n1277_;
  assign po155 = new_n1276_;
  assign po156 = new_n1275_;
  assign po157 = new_n1274_;
  assign po158 = new_n1273_;
  assign po159 = new_n1272_;
  assign po160 = new_n1271_;
  assign po161 = new_n1270_;
  assign po162 = new_n1269_;
  assign po163 = new_n1268_;
  assign po164 = new_n1267_;
  assign po165 = new_n1266_;
  assign po166 = new_n1265_;
  assign po167 = new_n1264_;
  assign po168 = new_n1263_;
  assign po169 = new_n1262_;
  assign po170 = new_n1261_;
  assign po171 = new_n1260_;
  assign po172 = new_n1259_;
  assign po173 = new_n1258_;
  assign po174 = new_n1257_;
  assign po175 = new_n1256_;
  assign po176 = new_n1255_;
  assign po177 = new_n1254_;
  assign po178 = new_n1253_;
  assign po179 = new_n1252_;
  assign po180 = new_n1251_;
  assign po181 = new_n1250_;
  assign po182 = new_n1249_;
  assign po183 = new_n1248_;
  assign po184 = new_n811_;
  assign po185 = new_n840_;
  assign po186 = new_n1375_;
  assign po187 = new_n1360_;
  assign po188 = new_n1334_;
  assign po189 = new_n1332_;
  assign po190 = new_n1338_;
  assign po191 = new_n1336_;
  assign po192 = new_n1342_;
  assign po193 = new_n1340_;
  assign po194 = new_n1346_;
  assign po195 = new_n1344_;
  assign po196 = new_n1350_;
  assign po197 = new_n1348_;
  assign po198 = new_n1356_;
  assign po199 = new_n1354_;
  assign po200 = new_n1357_;
  assign po201 = new_n1358_;
  assign po202 = new_n1361_;
  assign po203 = new_n1362_;
  assign po204 = new_n1363_;
  assign po205 = new_n1364_;
  assign po206 = new_n1365_;
  assign po207 = new_n1366_;
  assign po208 = new_n1367_;
  assign po209 = new_n1368_;
  assign po210 = new_n1369_;
  assign po211 = new_n1370_;
  assign po212 = new_n1371_;
  assign po213 = new_n1372_;
  assign po214 = new_n1373_;
  assign po215 = new_n1374_;
  assign po216 = new_n1287_;
  assign po217 = new_n1288_;
  assign po218 = new_n1289_;
  assign po219 = new_n1290_;
  assign po220 = new_n1291_;
  assign po221 = new_n1292_;
  assign po222 = new_n1293_;
  assign po223 = new_n1308_;
  assign po224 = new_n1295_;
  assign po225 = new_n1296_;
  assign po226 = new_n1297_;
  assign po227 = new_n1298_;
  assign po228 = new_n1299_;
  assign po229 = new_n1300_;
  assign po230 = new_n1301_;
  assign po231 = new_n1302_;
  assign po232 = new_n1303_;
  assign po233 = new_n1304_;
  assign po234 = new_n1305_;
  assign po235 = new_n1306_;
  assign po236 = new_n1314_;
  assign po237 = new_n1312_;
  assign po238 = new_n1320_;
  assign po239 = new_n1318_;
  assign po240 = new_n1326_;
  assign po241 = new_n1324_;
  assign po242 = new_n1330_;
  assign po243 = new_n1328_;
  assign po244 = new_n1286_;
  assign new_n747_ = new_n1395_ ? pi016 : (pi186 ^ new_n826_);
  assign new_n748_ = new_n1395_ ? pi007 : (pi187 ^ new_n828_);
  assign new_n749_ = new_n1395_ ? pi066 : (pi188 ^ new_n817_);
  assign new_n750_ = new_n1395_ ? (pi170 ^ new_n830_) : (~pi198 & pi067);
  assign new_n751_ = new_n1395_ ? (pi178 ^ new_n825_) : (~pi198 & pi069);
  assign new_n752_ = new_n1395_ ? (pi186 ^ new_n826_) : (~pi198 & pi071);
  assign new_n753_ = new_n1395_ ? (pi194 ^ new_n834_) : (~pi198 & pi073);
  assign new_n754_ = new_n1395_ ? (pi169 ^ new_n836_) : (pi198 ? pi067 : pi075);
  assign new_n755_ = new_n1395_ ? (pi177 ^ new_n838_) : (pi198 ? pi069 : pi077);
  assign new_n756_ = new_n1395_ ? (pi185 ^ new_n833_) : (pi198 ? pi071 : pi079);
  assign new_n757_ = new_n1395_ ? (pi193 ^ new_n837_) : (pi198 ? pi073 : pi081);
  assign new_n758_ = new_n1395_ ? (pi168 ^ new_n812_) : (pi198 ? pi075 : pi083);
  assign new_n759_ = new_n1395_ ? (pi176 ^ new_n820_) : (pi198 ? pi077 : pi085);
  assign new_n760_ = new_n1395_ ? (pi184 ^ new_n819_) : (pi198 ? pi079 : pi087);
  assign new_n761_ = new_n1395_ ? (pi192 ^ new_n831_) : (pi198 ? pi081 : pi089);
  assign new_n762_ = new_n1395_ ? (pi167 ^ new_n835_) : (pi198 ? pi083 : pi091);
  assign new_n763_ = new_n1395_ ? (pi175 ^ new_n832_) : (pi198 ? pi085 : pi093);
  assign new_n764_ = new_n1395_ ? (pi183 ^ new_n815_) : (pi198 ? pi087 : pi095);
  assign new_n765_ = new_n1395_ ? (pi191 ^ new_n842_) : (pi198 ? pi089 : pi097);
  assign new_n766_ = new_n1395_ ? (pi166 ^ new_n818_) : (pi198 ? pi091 : pi099);
  assign new_n767_ = new_n1395_ ? (pi174 ^ new_n814_) : (pi198 ? pi093 : pi101);
  assign new_n768_ = new_n1395_ ? (pi182 ^ new_n841_) : (pi198 ? pi095 : pi103);
  assign new_n769_ = new_n1395_ ? (pi190 ^ new_n839_) : (pi198 ? pi097 : pi105);
  assign new_n770_ = new_n1395_ ? (pi165 ^ new_n822_) : (pi198 ? pi099 : pi107);
  assign new_n771_ = new_n1395_ ? (pi173 ^ new_n816_) : (pi198 ? pi101 : pi109);
  assign new_n772_ = new_n1395_ ? (pi181 ^ new_n829_) : (pi198 ? pi103 : pi111);
  assign new_n773_ = new_n1395_ ? (pi189 ^ new_n821_) : (pi198 ? pi105 : pi113);
  assign new_n774_ = new_n1395_ ? (pi164 ^ new_n823_) : (pi198 ? pi107 : pi115);
  assign new_n775_ = new_n1395_ ? (pi172 ^ new_n824_) : (pi198 ? pi109 : pi117);
  assign new_n776_ = new_n1395_ ? (pi180 ^ new_n813_) : (pi198 ? pi111 : pi119);
  assign new_n777_ = new_n1395_ ? (pi188 ^ new_n817_) : (pi198 ? pi113 : pi121);
  assign new_n778_ = new_n1395_ ? (pi163 ^ new_n844_) : (pi198 ? pi115 : pi123);
  assign new_n779_ = new_n1395_ ? (pi171 ^ new_n843_) : (pi198 ? pi117 : pi125);
  assign new_n780_ = new_n1395_ ? (pi179 ^ new_n827_) : (pi198 ? pi119 : pi127);
  assign new_n781_ = new_n1395_ ? (pi187 ^ new_n828_) : (pi198 ? pi121 : pi129);
  assign new_n782_ = new_n1395_ ? pi001 : (pi163 ^ new_n844_);
  assign new_n783_ = new_n1395_ ? pi060 : (pi164 ^ new_n823_);
  assign new_n784_ = new_n1395_ ? pi052 : (pi165 ^ new_n822_);
  assign new_n785_ = new_n1395_ ? pi044 : (pi166 ^ new_n818_);
  assign new_n786_ = new_n1395_ ? pi036 : (pi167 ^ new_n835_);
  assign new_n787_ = new_n1395_ ? pi028 : (pi168 ^ new_n812_);
  assign new_n788_ = new_n1395_ ? pi020 : (pi169 ^ new_n836_);
  assign new_n789_ = new_n1395_ ? pi012 : (pi170 ^ new_n830_);
  assign new_n790_ = new_n1395_ ? pi003 : (pi171 ^ new_n843_);
  assign new_n791_ = new_n1395_ ? pi062 : (pi172 ^ new_n824_);
  assign new_n792_ = new_n1395_ ? pi054 : (pi173 ^ new_n816_);
  assign new_n793_ = new_n1395_ ? pi046 : (pi174 ^ new_n814_);
  assign new_n794_ = new_n1395_ ? pi038 : (pi175 ^ new_n832_);
  assign new_n795_ = new_n1395_ ? pi058 : (pi189 ^ new_n821_);
  assign new_n796_ = new_n1395_ ? pi050 : (pi190 ^ new_n839_);
  assign new_n797_ = new_n1395_ ? pi042 : (pi191 ^ new_n842_);
  assign new_n798_ = new_n1395_ ? pi034 : (pi192 ^ new_n831_);
  assign new_n799_ = new_n1395_ ? pi026 : (pi193 ^ new_n837_);
  assign new_n800_ = new_n1395_ ? pi018 : (pi194 ^ new_n834_);
  assign new_n801_ = new_n1395_ ? pi024 : (pi185 ^ new_n833_);
  assign new_n802_ = new_n1395_ ? pi032 : (pi184 ^ new_n819_);
  assign new_n803_ = new_n1395_ ? pi040 : (pi183 ^ new_n815_);
  assign new_n804_ = new_n1395_ ? pi048 : (pi182 ^ new_n841_);
  assign new_n805_ = new_n1395_ ? pi056 : (pi181 ^ new_n829_);
  assign new_n806_ = new_n1395_ ? pi064 : (pi180 ^ new_n813_);
  assign new_n807_ = new_n1395_ ? pi005 : (pi179 ^ new_n827_);
  assign new_n808_ = new_n1395_ ? pi014 : (pi178 ^ new_n825_);
  assign new_n809_ = new_n1395_ ? pi022 : (pi177 ^ new_n838_);
  assign new_n810_ = new_n1395_ ? pi030 : (pi176 ^ new_n820_);
  assign new_n811_ = ~new_n1407_ & ~pi008 & ((pi195 & (~pi196 | ~pi198 | ~pi197)) | (~pi195 & pi196 & pi198 & pi197));
  assign new_n812_ = (~new_n1422_ & (new_n1421_ ? (~new_n1425_ & (new_n1423_ ? (~new_n1424_ & new_n1426_) : (new_n1424_ & ~new_n1426_))) : (new_n1424_ & new_n1425_ & (~new_n1423_ ^ new_n1426_)))) | new_n1121_ | new_n1122_ | new_n1123_ | new_n1128_ | new_n1129_ | new_n1130_ | new_n1131_ | new_n1132_ | new_n1133_ | new_n1136_ | new_n1137_ | new_n1138_ | new_n1139_ | new_n1141_ | new_n1143_ | new_n1146_ | new_n1147_ | new_n1148_ | new_n1150_ | new_n1151_ | new_n1153_ | new_n1154_ | new_n1155_ | new_n1157_ | new_n1158_ | new_n1159_ | new_n1162_ | new_n1163_;
  assign new_n813_ = (~new_n1422_ & ((new_n1421_ & ((~new_n1423_ & ~new_n1424_ & ~new_n1425_ & new_n1426_) | (new_n1423_ & new_n1424_ & new_n1425_ & ~new_n1426_))) | (~new_n1421_ & ~new_n1423_ & ~new_n1424_ & new_n1425_ & ~new_n1426_))) | new_n1122_ | new_n1123_ | new_n1124_ | new_n1125_ | new_n1127_ | new_n1128_ | new_n1131_ | new_n1132_ | new_n1134_ | new_n1135_ | new_n1136_ | new_n1139_ | new_n1140_ | new_n1141_ | new_n1143_ | new_n1144_ | new_n1147_ | new_n1148_ | new_n1149_ | new_n1151_ | new_n1152_ | new_n1154_ | new_n1155_ | new_n1156_ | new_n1158_ | new_n1161_ | new_n1163_ | new_n1164_ | (~new_n1421_ & new_n1422_ & new_n1423_ & new_n1424_ & new_n1425_ & new_n1426_);
  assign new_n814_ = new_n1121_ | new_n1123_ | new_n1124_ | new_n1126_ | new_n1127_ | new_n1129_ | new_n1131_ | new_n1132_ | new_n1133_ | new_n1135_ | new_n1136_ | new_n1138_ | new_n1140_ | new_n1142_ | new_n1143_ | new_n1144_ | new_n1145_ | new_n1150_ | new_n1151_ | new_n1152_ | new_n1153_ | new_n1155_ | new_n1157_ | new_n1158_ | new_n1160_ | new_n1161_ | new_n1162_ | new_n1164_ | (~new_n1422_ & ((~new_n1423_ & ((new_n1421_ & new_n1425_ & (new_n1424_ ^ new_n1426_)) | (~new_n1425_ & new_n1426_ & ~new_n1421_ & ~new_n1424_))) | (~new_n1421_ & new_n1423_ & new_n1424_ & new_n1425_ & ~new_n1426_)));
  assign new_n815_ = new_n1074_ | new_n1075_ | new_n1076_ | new_n1078_ | new_n1080_ | new_n1081_ | new_n1083_ | new_n1084_ | new_n1086_ | new_n1089_ | new_n1091_ | new_n1092_ | new_n1093_ | new_n1094_ | new_n1096_ | new_n1097_ | new_n1099_ | new_n1100_ | new_n1102_ | new_n1103_ | new_n1104_ | new_n1106_ | new_n1108_ | new_n1110_ | new_n1112_ | new_n1113_ | new_n1114_ | new_n1116_ | (~new_n1416_ & ~new_n1418_ & (~new_n1417_ ^ new_n1420_) & (~new_n1415_ ^ new_n1419_));
  assign new_n816_ = (new_n1416_ & new_n1417_ & ((new_n1415_ & new_n1419_ & (new_n1418_ ^ new_n1420_)) | (~new_n1419_ & new_n1420_ & ~new_n1415_ & ~new_n1418_))) | new_n1073_ | new_n1074_ | new_n1075_ | new_n1077_ | new_n1080_ | new_n1082_ | new_n1083_ | new_n1085_ | new_n1086_ | new_n1088_ | new_n1089_ | new_n1090_ | new_n1093_ | new_n1094_ | new_n1095_ | new_n1098_ | new_n1099_ | new_n1100_ | new_n1101_ | new_n1102_ | new_n1103_ | new_n1106_ | new_n1107_ | new_n1109_ | new_n1110_ | new_n1113_ | new_n1114_ | new_n1115_ | (~new_n1415_ & ~new_n1416_ & ~new_n1417_ & new_n1418_ & ~new_n1419_ & ~new_n1420_);
  assign new_n817_ = (~new_n1416_ & ~new_n1419_ & ((new_n1415_ & ~new_n1418_ & (~new_n1417_ ^ new_n1420_)) | (~new_n1415_ & new_n1417_ & new_n1418_ & new_n1420_))) | new_n1073_ | new_n1075_ | new_n1076_ | new_n1077_ | new_n1079_ | new_n1080_ | new_n1081_ | new_n1084_ | new_n1085_ | new_n1086_ | new_n1087_ | new_n1090_ | new_n1091_ | new_n1093_ | new_n1095_ | new_n1096_ | new_n1098_ | new_n1099_ | new_n1102_ | new_n1104_ | new_n1105_ | new_n1107_ | new_n1108_ | new_n1110_ | new_n1111_ | new_n1112_ | new_n1113_ | new_n1115_ | (~new_n1415_ & new_n1416_ & new_n1417_ & new_n1418_ & new_n1419_ & ~new_n1420_);
  assign new_n818_ = new_n1024_ | new_n1026_ | new_n1028_ | new_n1283_ | new_n1031_ | new_n1032_ | new_n1033_ | new_n1036_ | new_n1037_ | new_n1038_ | new_n1040_ | new_n1041_ | new_n1042_ | new_n1043_ | new_n1047_ | new_n1048_ | new_n1049_ | new_n1050_ | new_n1052_ | new_n1054_ | new_n1056_ | new_n1058_ | new_n1060_ | new_n1061_ | new_n1064_ | new_n1066_ | new_n1067_ | new_n1068_ | (~new_n1392_ & ((~new_n1393_ & ((new_n1412_ & (new_n1391_ ? (new_n1414_ & ~new_n1394_) : (~new_n1414_ & new_n1394_))) | (new_n1414_ & new_n1394_ & ~new_n1412_ & ~new_n1391_))) | (new_n1414_ & new_n1393_ & ~new_n1394_ & ~new_n1412_ & new_n1391_)));
  assign new_n819_ = new_n1025_ | new_n1026_ | new_n1028_ | new_n1030_ | new_n1031_ | new_n1032_ | new_n1034_ | new_n1035_ | new_n1036_ | new_n1037_ | new_n1041_ | new_n1043_ | new_n1044_ | new_n1045_ | new_n1047_ | new_n1048_ | new_n1051_ | new_n1052_ | new_n1053_ | new_n1055_ | new_n1056_ | new_n1057_ | new_n1061_ | new_n1062_ | new_n1063_ | new_n1064_ | new_n1066_ | new_n1067_ | (~new_n1391_ & (new_n1392_ ? (~new_n1414_ & ~new_n1394_) : (new_n1414_ & new_n1394_)) & (new_n1412_ ^ new_n1393_));
  assign new_n820_ = (new_n1391_ & ((new_n1412_ & ~new_n1393_ & (new_n1392_ ? (~new_n1414_ & ~new_n1394_) : (new_n1414_ & new_n1394_))) | (~new_n1412_ & ~new_n1392_ & ~new_n1414_ & new_n1393_ & new_n1394_))) | new_n1026_ | new_n1027_ | new_n1283_ | new_n1030_ | new_n1032_ | new_n1033_ | new_n1034_ | new_n1036_ | new_n1037_ | new_n1039_ | new_n1040_ | new_n1042_ | new_n1044_ | new_n1045_ | new_n1046_ | new_n1048_ | new_n1049_ | new_n1051_ | new_n1052_ | new_n1054_ | new_n1055_ | new_n1057_ | new_n1059_ | new_n1060_ | new_n1061_ | new_n1063_ | new_n1066_ | new_n1068_ | (~new_n1414_ & new_n1393_ & ~new_n1394_ & ~new_n1412_ & ~new_n1391_ & ~new_n1392_);
  assign new_n821_ = new_n881_ | new_n914_ | new_n885_ | new_n886_ | new_n887_ | new_n889_ | new_n890_ | new_n891_ | new_n892_ | new_n930_ | new_n893_ | new_n896_ | new_n899_ | new_n900_ | new_n901_ | new_n904_ | new_n906_ | new_n907_ | new_n908_ | new_n910_ | new_n913_ | new_n915_ | new_n917_ | new_n918_ | new_n919_ | new_n921_ | new_n922_ | new_n923_ | (~new_n1378_ & new_n1376_ & new_n1382_ & new_n1400_ & new_n1383_ & new_n1401_) | (~new_n1382_ & ~new_n1400_ & ((new_n1378_ & (new_n1376_ ? (new_n1383_ & ~new_n1401_) : (~new_n1383_ & new_n1401_))) | (~new_n1383_ & ~new_n1401_ & ~new_n1378_ & new_n1376_)));
  assign new_n822_ = new_n880_ | new_n882_ | new_n920_ | new_n914_ | new_n885_ | new_n889_ | new_n890_ | new_n892_ | new_n893_ | new_n894_ | new_n895_ | new_n897_ | new_n899_ | new_n900_ | new_n902_ | new_n906_ | new_n907_ | new_n908_ | new_n911_ | new_n912_ | new_n913_ | new_n976_ | new_n916_ | new_n918_ | new_n919_ | new_n994_ | new_n921_ | new_n922_ | (new_n1376_ & ~new_n1383_ & ((new_n1400_ & (new_n1378_ ? (~new_n1382_ ^ new_n1401_) : (new_n1382_ & ~new_n1401_))) | (~new_n1400_ & new_n1401_ & ~new_n1378_ & ~new_n1382_)));
  assign new_n823_ = new_n1005_ | new_n973_ | new_n925_ | new_n877_ | new_n927_ | new_n1188_ | new_n1184_ | new_n1183_ | new_n1182_ | new_n1281_ | new_n1181_ | new_n1179_ | new_n1177_ | new_n1176_ | new_n1174_ | new_n1173_ | new_n1172_ | new_n1170_ | new_n1169_ | new_n1166_ | new_n1165_ | new_n1120_ | new_n1119_ | new_n1118_ | new_n1280_ | new_n926_ | new_n1191_ | new_n1117_ | (~new_n1381_ & (new_n1397_ ? ((~new_n1409_ & new_n1411_ & new_n1380_ & new_n1398_) | (~new_n1380_ & ~new_n1398_ & new_n1409_ & ~new_n1411_)) : (new_n1398_ & new_n1409_ & (~new_n1380_ ^ new_n1411_))));
  assign new_n824_ = new_n1282_ | new_n1065_ | new_n925_ | new_n877_ | new_n927_ | new_n1189_ | new_n1187_ | new_n1186_ | new_n1184_ | new_n1181_ | new_n1180_ | new_n1178_ | new_n1177_ | new_n1176_ | new_n1173_ | new_n1172_ | new_n1171_ | new_n1169_ | new_n1165_ | new_n1119_ | new_n1118_ | new_n1072_ | new_n1280_ | new_n1071_ | new_n1070_ | new_n1191_ | new_n1117_ | new_n1069_ | (~new_n1381_ & (new_n1397_ ? (new_n1398_ & (new_n1380_ ? (~new_n1409_ & ~new_n1411_) : (new_n1409_ & new_n1411_))) : (new_n1380_ & ~new_n1398_ & (~new_n1409_ ^ new_n1411_))));
  assign new_n825_ = new_n1282_ | new_n1065_ | new_n1020_ | new_n1005_ | new_n925_ | new_n877_ | new_n927_ | new_n1189_ | new_n1188_ | new_n1186_ | new_n1185_ | new_n1182_ | new_n1281_ | new_n1180_ | new_n1179_ | new_n1178_ | new_n1176_ | new_n1175_ | new_n1173_ | new_n1170_ | new_n1169_ | new_n1168_ | new_n1165_ | new_n1120_ | new_n1072_ | new_n1280_ | new_n1070_ | new_n926_ | (~new_n1381_ & ((~new_n1398_ & ((new_n1397_ & ~new_n1409_ & (~new_n1380_ ^ new_n1411_)) | (new_n1409_ & ~new_n1411_ & ~new_n1397_ & ~new_n1380_))) | (~new_n1397_ & ~new_n1380_ & new_n1398_ & new_n1409_ & new_n1411_)));
  assign new_n826_ = new_n1282_ | new_n1020_ | new_n973_ | new_n877_ | new_n1189_ | new_n1188_ | new_n1187_ | new_n1185_ | new_n1184_ | new_n1183_ | new_n1281_ | new_n1180_ | new_n1179_ | new_n1177_ | new_n1176_ | new_n1175_ | new_n1174_ | new_n1171_ | new_n1169_ | new_n1168_ | new_n1166_ | new_n1119_ | new_n1072_ | new_n1280_ | new_n1071_ | new_n926_ | new_n1191_ | new_n1069_ | (new_n1398_ & ((~new_n1381_ & ((new_n1397_ & ~new_n1380_ & (new_n1409_ ^ new_n1411_)) | (new_n1409_ & ~new_n1411_ & ~new_n1397_ & new_n1380_))) | (~new_n1397_ & new_n1381_ & new_n1380_ & new_n1409_ & new_n1411_)));
  assign new_n827_ = (new_n1378_ & ~new_n1382_ & ~new_n1383_ & (new_n1376_ ? (~new_n1400_ & new_n1401_) : (new_n1400_ & ~new_n1401_))) | new_n882_ | new_n920_ | new_n885_ | new_n886_ | new_n887_ | new_n888_ | new_n889_ | new_n891_ | new_n892_ | new_n894_ | new_n896_ | new_n897_ | new_n898_ | new_n900_ | new_n901_ | new_n902_ | new_n906_ | new_n909_ | new_n910_ | new_n912_ | new_n913_ | new_n915_ | new_n916_ | new_n918_ | new_n919_ | new_n994_ | new_n923_ | new_n924_ | (~new_n1378_ & new_n1382_ & ~new_n1400_ & new_n1383_ & (new_n1376_ ^ new_n1401_));
  assign new_n828_ = (new_n1387_ & ~new_n1408_ & new_n1389_ & (new_n1388_ ? (new_n1410_ & ~new_n1390_) : (~new_n1410_ & new_n1390_))) | new_n977_ | new_n979_ | new_n980_ | new_n984_ | new_n985_ | new_n986_ | new_n987_ | new_n988_ | new_n989_ | new_n990_ | new_n992_ | new_n1190_ | new_n995_ | new_n997_ | new_n999_ | new_n1000_ | new_n1001_ | new_n1003_ | new_n1004_ | new_n1167_ | new_n1008_ | new_n1009_ | new_n1010_ | new_n1012_ | new_n1013_ | new_n1015_ | new_n1016_ | new_n1017_ | (~new_n1387_ & new_n1408_ & ~new_n1389_ & (new_n1388_ ? (new_n1410_ & new_n1390_) : (~new_n1410_ & ~new_n1390_)));
  assign new_n829_ = new_n977_ | new_n978_ | new_n981_ | new_n982_ | new_n984_ | new_n985_ | new_n986_ | new_n988_ | new_n990_ | new_n991_ | new_n992_ | new_n993_ | new_n1190_ | new_n998_ | new_n1001_ | new_n1002_ | new_n1003_ | new_n1167_ | new_n1284_ | new_n1006_ | new_n1008_ | new_n1010_ | new_n1011_ | new_n1012_ | new_n1013_ | new_n1014_ | new_n1015_ | new_n1018_ | (~new_n1387_ & ~new_n1408_ & ~new_n1388_ & new_n1410_ & ~new_n1389_ & ~new_n1390_) | (~new_n1410_ & ((new_n1387_ & ((new_n1408_ & new_n1388_ & new_n1389_ & new_n1390_) | (~new_n1408_ & ~new_n1388_ & ~new_n1389_ & ~new_n1390_))) | (~new_n1387_ & ~new_n1408_ & new_n1388_ & ~new_n1389_ & new_n1390_)));
  assign new_n830_ = new_n978_ | new_n979_ | new_n980_ | new_n981_ | new_n983_ | new_n984_ | new_n986_ | new_n988_ | new_n989_ | new_n991_ | new_n1190_ | new_n995_ | new_n996_ | new_n998_ | new_n999_ | new_n1000_ | new_n1002_ | new_n1003_ | new_n1006_ | new_n1007_ | new_n1008_ | new_n1009_ | new_n1011_ | new_n1012_ | new_n1014_ | new_n1015_ | new_n1017_ | new_n1019_ | (~new_n1408_ & (new_n1387_ ? ((~new_n1389_ & new_n1390_ & new_n1388_ & new_n1410_) | (~new_n1388_ & ~new_n1410_ & new_n1389_ & ~new_n1390_)) : (~new_n1388_ & ~new_n1389_ & (~new_n1410_ ^ new_n1390_))));
  assign new_n831_ = (~new_n1408_ & (new_n1387_ ? (~new_n1389_ & (new_n1388_ ? (~new_n1410_ & new_n1390_) : (new_n1410_ & ~new_n1390_))) : (new_n1410_ & new_n1389_ & (~new_n1388_ ^ new_n1390_)))) | new_n978_ | new_n980_ | new_n982_ | new_n983_ | new_n984_ | new_n985_ | new_n987_ | new_n989_ | new_n991_ | new_n992_ | new_n993_ | new_n1190_ | new_n996_ | new_n997_ | new_n999_ | new_n1001_ | new_n1002_ | new_n1003_ | new_n1004_ | new_n1284_ | new_n1007_ | new_n1009_ | new_n1011_ | new_n1013_ | new_n1015_ | new_n1016_ | new_n1018_ | new_n1019_;
  assign new_n832_ = new_n1023_ | new_n931_ | new_n932_ | new_n934_ | new_n937_ | new_n939_ | new_n940_ | new_n941_ | new_n943_ | new_n944_ | new_n945_ | new_n947_ | new_n948_ | new_n949_ | new_n952_ | new_n954_ | new_n956_ | new_n957_ | new_n958_ | new_n960_ | new_n961_ | new_n963_ | new_n964_ | new_n966_ | new_n968_ | new_n970_ | new_n971_ | new_n972_ | (new_n1402_ & (~new_n1384_ ^ new_n1386_) & (new_n1385_ ? (new_n1404_ & ~new_n1406_) : (~new_n1404_ & new_n1406_)));
  assign new_n833_ = new_n1023_ | new_n932_ | new_n933_ | new_n934_ | new_n936_ | new_n938_ | new_n940_ | new_n942_ | new_n944_ | new_n945_ | new_n946_ | new_n947_ | new_n1029_ | new_n949_ | new_n951_ | new_n952_ | new_n955_ | new_n956_ | new_n958_ | new_n959_ | new_n960_ | new_n962_ | new_n963_ | new_n964_ | new_n965_ | new_n969_ | new_n971_ | new_n972_ | (new_n1402_ & (new_n1404_ ? (~new_n1386_ & new_n1406_) : (new_n1386_ & ~new_n1406_)) & (new_n1384_ ^ ~new_n1385_));
  assign new_n834_ = new_n1023_ | new_n931_ | new_n933_ | new_n935_ | new_n937_ | new_n938_ | new_n940_ | new_n941_ | new_n942_ | new_n943_ | new_n945_ | new_n946_ | new_n947_ | new_n950_ | new_n953_ | new_n955_ | new_n956_ | new_n957_ | new_n958_ | new_n959_ | new_n961_ | new_n962_ | new_n963_ | new_n966_ | new_n967_ | new_n968_ | new_n969_ | new_n971_ | (~new_n1404_ & (new_n1384_ ? (new_n1386_ & (new_n1402_ ? (~new_n1385_ & ~new_n1406_) : (new_n1385_ & new_n1406_))) : (new_n1402_ & ~new_n1386_ & (~new_n1385_ ^ new_n1406_))));
  assign new_n835_ = new_n871_ | new_n859_ | new_n879_ | new_n862_ | new_n865_ | new_n884_ | new_n869_ | new_n872_ | new_n873_ | new_n874_ | new_n875_ | new_n876_ | new_n928_ | new_n1022_ | new_n1021_ | new_n883_ | new_n878_ | new_n870_ | new_n860_ | new_n849_ | new_n845_ | new_n846_ | new_n852_ | new_n848_ | new_n857_ | new_n853_ | new_n854_ | new_n855_ | (~new_n1427_ & ((new_n1379_ & ((new_n1377_ & ~new_n1399_ & (~new_n1413_ ^ ~new_n1396_)) | (new_n1413_ & new_n1396_ & ~new_n1377_ & new_n1399_))) | (~new_n1377_ & new_n1399_ & ~new_n1413_ & ~new_n1379_ & new_n1396_)));
  assign new_n836_ = (new_n1404_ & ((new_n1384_ & new_n1385_ & (new_n1402_ ? (~new_n1386_ & ~new_n1406_) : (new_n1386_ & new_n1406_))) | (~new_n1384_ & new_n1402_ & ~new_n1385_ & ~new_n1386_ & ~new_n1406_))) | new_n931_ | new_n932_ | new_n935_ | new_n936_ | new_n938_ | new_n939_ | new_n940_ | new_n941_ | new_n942_ | new_n945_ | new_n948_ | new_n1029_ | new_n949_ | new_n950_ | new_n951_ | new_n953_ | new_n954_ | new_n955_ | new_n957_ | new_n958_ | new_n960_ | new_n963_ | new_n965_ | new_n966_ | new_n967_ | new_n969_ | new_n970_ | new_n972_ | (~new_n1384_ & ~new_n1402_ & ~new_n1385_ & ~new_n1404_ & new_n1386_ & new_n1406_);
  assign new_n837_ = (new_n1379_ & ((new_n1377_ & new_n1399_ & ~new_n1427_ & (~new_n1413_ ^ new_n1396_)) | (~new_n1377_ & ~new_n1399_ & new_n1413_ & new_n1427_ & new_n1396_))) | new_n866_ | new_n856_ | new_n862_ | new_n864_ | new_n865_ | new_n867_ | new_n868_ | new_n869_ | new_n903_ | new_n872_ | new_n873_ | new_n876_ | new_n928_ | new_n1022_ | new_n1021_ | new_n975_ | new_n974_ | new_n883_ | new_n847_ | new_n850_ | new_n845_ | new_n846_ | new_n852_ | new_n858_ | new_n857_ | new_n861_ | new_n854_ | new_n855_ | (~new_n1377_ & ~new_n1399_ & ~new_n1413_ & new_n1427_ & ~new_n1379_ & new_n1396_);
  assign new_n838_ = (~new_n1379_ & ((new_n1377_ & ~new_n1427_ & (new_n1399_ ? (new_n1413_ & new_n1396_) : (~new_n1413_ & ~new_n1396_))) | (~new_n1377_ & new_n1399_ & ~new_n1413_ & new_n1427_ & new_n1396_))) | new_n866_ | new_n871_ | new_n859_ | new_n863_ | new_n864_ | new_n865_ | new_n884_ | new_n868_ | new_n869_ | new_n903_ | new_n873_ | new_n875_ | new_n905_ | new_n928_ | new_n975_ | new_n974_ | new_n929_ | new_n883_ | new_n878_ | new_n860_ | new_n850_ | new_n849_ | new_n845_ | new_n846_ | new_n851_ | new_n861_ | new_n853_ | new_n855_ | (~new_n1427_ & new_n1379_ & new_n1396_ & new_n1377_ & ~new_n1399_ & new_n1413_);
  assign new_n839_ = new_n1121_ | new_n1123_ | new_n1124_ | new_n1125_ | new_n1126_ | new_n1128_ | new_n1130_ | new_n1132_ | new_n1133_ | new_n1134_ | new_n1137_ | new_n1140_ | new_n1141_ | new_n1142_ | new_n1144_ | new_n1145_ | new_n1146_ | new_n1147_ | new_n1149_ | new_n1150_ | new_n1151_ | new_n1154_ | new_n1156_ | new_n1157_ | new_n1158_ | new_n1159_ | new_n1160_ | new_n1164_ | (new_n1424_ & (new_n1421_ ? (new_n1423_ & (new_n1422_ ? (new_n1425_ & ~new_n1426_) : (~new_n1425_ & new_n1426_))) : (~new_n1422_ & ~new_n1423_ & (~new_n1425_ ^ new_n1426_))));
  assign new_n840_ = ~new_n1407_ & ~pi008 & (~pi196 ^ (~pi198 | ~pi197));
  assign new_n841_ = (~new_n1379_ & ((new_n1377_ & new_n1413_ & ~new_n1396_ & (new_n1399_ ^ new_n1427_)) | (~new_n1377_ & ~new_n1399_ & ~new_n1413_ & ~new_n1427_ & new_n1396_))) | new_n866_ | new_n856_ | new_n871_ | new_n879_ | new_n863_ | new_n865_ | new_n884_ | new_n867_ | new_n869_ | new_n903_ | new_n874_ | new_n876_ | new_n905_ | new_n928_ | new_n1022_ | new_n975_ | new_n929_ | new_n878_ | new_n870_ | new_n847_ | new_n849_ | new_n846_ | new_n852_ | new_n848_ | new_n858_ | new_n851_ | new_n861_ | new_n854_ | (~new_n1427_ & new_n1379_ & new_n1396_ & ~new_n1377_ & new_n1399_ & ~new_n1413_);
  assign new_n842_ = new_n1024_ | new_n1025_ | new_n1026_ | new_n1027_ | new_n1283_ | new_n1031_ | new_n1034_ | new_n1035_ | new_n1036_ | new_n1038_ | new_n1039_ | new_n1042_ | new_n1043_ | new_n1044_ | new_n1046_ | new_n1047_ | new_n1048_ | new_n1050_ | new_n1053_ | new_n1054_ | new_n1055_ | new_n1058_ | new_n1059_ | new_n1061_ | new_n1062_ | new_n1063_ | new_n1064_ | new_n1068_ | (new_n1392_ & (new_n1412_ ? ((~new_n1393_ & new_n1394_ & new_n1391_ & new_n1414_) | (new_n1393_ & ~new_n1394_ & ~new_n1391_ & ~new_n1414_)) : (new_n1414_ & new_n1393_ & (~new_n1391_ ^ new_n1394_))));
  assign new_n843_ = new_n880_ | new_n881_ | new_n882_ | new_n885_ | new_n887_ | new_n888_ | new_n890_ | new_n891_ | new_n930_ | new_n895_ | new_n897_ | new_n898_ | new_n899_ | new_n900_ | new_n901_ | new_n904_ | new_n906_ | new_n908_ | new_n909_ | new_n911_ | new_n912_ | new_n976_ | new_n915_ | new_n917_ | new_n919_ | new_n994_ | new_n922_ | new_n924_ | (~new_n1400_ & new_n1383_ & new_n1401_ & ~new_n1378_ & new_n1376_ & ~new_n1382_) | (new_n1382_ & ((new_n1400_ & new_n1383_ & ~new_n1401_ & ~new_n1378_ & new_n1376_) | (new_n1378_ & ~new_n1376_ & ~new_n1383_ & (~new_n1400_ ^ new_n1401_))));
  assign new_n844_ = new_n1073_ | new_n1074_ | new_n1075_ | new_n1076_ | new_n1078_ | new_n1079_ | new_n1082_ | new_n1084_ | new_n1085_ | new_n1087_ | new_n1088_ | new_n1089_ | new_n1092_ | new_n1093_ | new_n1095_ | new_n1096_ | new_n1097_ | new_n1100_ | new_n1101_ | new_n1102_ | new_n1105_ | new_n1107_ | new_n1108_ | new_n1109_ | new_n1111_ | new_n1113_ | new_n1114_ | new_n1116_ | (new_n1418_ & (new_n1415_ ? (~new_n1417_ & new_n1419_ & (new_n1416_ ^ new_n1420_)) : (new_n1417_ & ~new_n1419_ & (~new_n1416_ ^ new_n1420_))));
  assign new_n845_ = new_n1396_ & ~new_n1379_ & ~new_n1427_ & ~new_n1413_ & new_n1377_ & new_n1399_;
  assign new_n846_ = ~new_n1396_ & new_n1379_ & ~new_n1427_ & ~new_n1413_ & ~new_n1377_ & new_n1399_;
  assign new_n847_ = new_n1396_ & new_n1379_ & new_n1427_ & ~new_n1413_ & new_n1377_ & ~new_n1399_;
  assign new_n848_ = ~new_n1396_ & ~new_n1379_ & new_n1427_ & ~new_n1413_ & ~new_n1377_ & new_n1399_;
  assign new_n849_ = ~new_n1396_ & ~new_n1379_ & ~new_n1427_ & ~new_n1413_ & new_n1377_ & new_n1399_;
  assign new_n850_ = ~new_n1396_ & ~new_n1379_ & ~new_n1427_ & ~new_n1413_ & ~new_n1377_ & new_n1399_;
  assign new_n851_ = ~new_n1396_ & new_n1379_ & new_n1427_ & ~new_n1413_ & new_n1377_ & new_n1399_;
  assign new_n852_ = new_n1396_ & new_n1379_ & ~new_n1427_ & ~new_n1413_ & new_n1377_ & new_n1399_;
  assign new_n853_ = new_n1396_ & new_n1379_ & new_n1427_ & ~new_n1413_ & new_n1377_ & new_n1399_;
  assign new_n854_ = ~new_n1396_ & ~new_n1379_ & ~new_n1427_ & new_n1413_ & new_n1377_ & ~new_n1399_;
  assign new_n855_ = new_n1396_ & ~new_n1379_ & ~new_n1427_ & new_n1413_ & ~new_n1377_ & ~new_n1399_;
  assign new_n856_ = ~new_n1396_ & new_n1379_ & ~new_n1427_ & new_n1413_ & ~new_n1377_ & ~new_n1399_;
  assign new_n857_ = ~new_n1396_ & new_n1379_ & new_n1427_ & ~new_n1413_ & ~new_n1377_ & new_n1399_;
  assign new_n858_ = new_n1396_ & ~new_n1379_ & new_n1427_ & ~new_n1413_ & new_n1377_ & new_n1399_;
  assign new_n859_ = ~new_n1396_ & ~new_n1379_ & new_n1427_ & new_n1413_ & ~new_n1377_ & ~new_n1399_;
  assign new_n860_ = new_n1396_ & new_n1379_ & new_n1427_ & ~new_n1413_ & ~new_n1377_ & ~new_n1399_;
  assign new_n861_ = new_n1396_ & new_n1379_ & new_n1427_ & ~new_n1413_ & ~new_n1377_ & new_n1399_;
  assign new_n862_ = new_n1396_ & ~new_n1379_ & new_n1427_ & new_n1413_ & new_n1377_ & ~new_n1399_;
  assign new_n863_ = ~new_n1396_ & new_n1379_ & new_n1427_ & new_n1413_ & ~new_n1377_ & ~new_n1399_;
  assign new_n864_ = ~new_n1396_ & new_n1379_ & new_n1427_ & new_n1413_ & new_n1377_ & ~new_n1399_;
  assign new_n865_ = new_n1396_ & new_n1379_ & new_n1427_ & new_n1413_ & new_n1377_ & ~new_n1399_;
  assign new_n866_ = new_n1396_ & ~new_n1379_ & ~new_n1427_ & new_n1413_ & new_n1377_ & ~new_n1399_;
  assign new_n867_ = new_n1396_ & ~new_n1379_ & ~new_n1427_ & new_n1413_ & ~new_n1377_ & new_n1399_;
  assign new_n868_ = ~new_n1396_ & new_n1379_ & ~new_n1427_ & new_n1413_ & ~new_n1377_ & new_n1399_;
  assign new_n869_ = ~new_n1396_ & new_n1379_ & ~new_n1427_ & new_n1413_ & new_n1377_ & new_n1399_;
  assign new_n870_ = ~new_n1396_ & new_n1379_ & new_n1427_ & ~new_n1413_ & ~new_n1377_ & ~new_n1399_;
  assign new_n871_ = new_n1396_ & new_n1379_ & ~new_n1427_ & new_n1413_ & ~new_n1377_ & ~new_n1399_;
  assign new_n872_ = ~new_n1396_ & ~new_n1379_ & new_n1427_ & new_n1413_ & new_n1377_ & new_n1399_;
  assign new_n873_ = new_n1396_ & ~new_n1379_ & new_n1427_ & new_n1413_ & ~new_n1377_ & new_n1399_;
  assign new_n874_ = new_n1396_ & ~new_n1379_ & new_n1427_ & new_n1413_ & new_n1377_ & new_n1399_;
  assign new_n875_ = ~new_n1396_ & new_n1379_ & new_n1427_ & new_n1413_ & new_n1377_ & new_n1399_;
  assign new_n876_ = new_n1396_ & new_n1379_ & new_n1427_ & new_n1413_ & ~new_n1377_ & new_n1399_;
  assign new_n877_ = new_n1411_ & new_n1409_ & ~new_n1398_ & ~new_n1380_ & ~new_n1397_ & ~new_n1381_;
  assign new_n878_ = new_n1396_ & ~new_n1379_ & new_n1427_ & ~new_n1413_ & new_n1377_ & ~new_n1399_;
  assign new_n879_ = new_n1396_ & ~new_n1379_ & new_n1427_ & new_n1413_ & ~new_n1377_ & ~new_n1399_;
  assign new_n880_ = ~new_n1401_ & ~new_n1383_ & ~new_n1400_ & ~new_n1382_ & ~new_n1378_ & ~new_n1376_;
  assign new_n881_ = ~new_n1401_ & ~new_n1383_ & new_n1400_ & ~new_n1382_ & ~new_n1378_ & ~new_n1376_;
  assign new_n882_ = ~new_n1401_ & new_n1383_ & new_n1400_ & ~new_n1382_ & ~new_n1378_ & ~new_n1376_;
  assign new_n883_ = ~new_n1396_ & ~new_n1379_ & new_n1427_ & ~new_n1413_ & new_n1377_ & ~new_n1399_;
  assign new_n884_ = ~new_n1396_ & ~new_n1379_ & ~new_n1427_ & new_n1413_ & ~new_n1377_ & new_n1399_;
  assign new_n885_ = ~new_n1401_ & ~new_n1383_ & new_n1400_ & new_n1382_ & ~new_n1378_ & ~new_n1376_;
  assign new_n886_ = ~new_n1401_ & new_n1383_ & new_n1400_ & new_n1382_ & ~new_n1378_ & ~new_n1376_;
  assign new_n887_ = ~new_n1401_ & new_n1383_ & ~new_n1400_ & ~new_n1382_ & ~new_n1378_ & new_n1376_;
  assign new_n888_ = ~new_n1401_ & ~new_n1383_ & new_n1400_ & ~new_n1382_ & ~new_n1378_ & new_n1376_;
  assign new_n889_ = ~new_n1401_ & new_n1383_ & new_n1400_ & ~new_n1382_ & ~new_n1378_ & new_n1376_;
  assign new_n890_ = ~new_n1401_ & ~new_n1383_ & ~new_n1400_ & new_n1382_ & ~new_n1378_ & new_n1376_;
  assign new_n891_ = new_n1401_ & ~new_n1383_ & ~new_n1400_ & ~new_n1382_ & ~new_n1378_ & ~new_n1376_;
  assign new_n892_ = new_n1401_ & new_n1383_ & ~new_n1400_ & ~new_n1382_ & ~new_n1378_ & ~new_n1376_;
  assign new_n893_ = new_n1401_ & ~new_n1383_ & ~new_n1400_ & new_n1382_ & ~new_n1378_ & ~new_n1376_;
  assign new_n894_ = new_n1401_ & ~new_n1383_ & new_n1400_ & new_n1382_ & ~new_n1378_ & ~new_n1376_;
  assign new_n895_ = new_n1401_ & new_n1383_ & new_n1400_ & new_n1382_ & ~new_n1378_ & ~new_n1376_;
  assign new_n896_ = new_n1401_ & ~new_n1383_ & new_n1400_ & ~new_n1382_ & ~new_n1378_ & new_n1376_;
  assign new_n897_ = new_n1401_ & new_n1383_ & new_n1400_ & ~new_n1382_ & ~new_n1378_ & new_n1376_;
  assign new_n898_ = new_n1401_ & ~new_n1383_ & ~new_n1400_ & new_n1382_ & ~new_n1378_ & new_n1376_;
  assign new_n899_ = new_n1401_ & new_n1383_ & ~new_n1400_ & new_n1382_ & ~new_n1378_ & new_n1376_;
  assign new_n900_ = new_n1401_ & ~new_n1383_ & new_n1400_ & new_n1382_ & ~new_n1378_ & new_n1376_;
  assign new_n901_ = ~new_n1401_ & ~new_n1383_ & ~new_n1400_ & ~new_n1382_ & new_n1378_ & ~new_n1376_;
  assign new_n902_ = ~new_n1401_ & new_n1383_ & ~new_n1400_ & ~new_n1382_ & new_n1378_ & ~new_n1376_;
  assign new_n903_ = ~new_n1396_ & ~new_n1379_ & new_n1427_ & new_n1413_ & ~new_n1377_ & new_n1399_;
  assign new_n904_ = ~new_n1401_ & new_n1383_ & new_n1400_ & ~new_n1382_ & new_n1378_ & ~new_n1376_;
  assign new_n905_ = new_n1396_ & new_n1379_ & new_n1427_ & new_n1413_ & new_n1377_ & new_n1399_;
  assign new_n906_ = ~new_n1401_ & new_n1383_ & ~new_n1400_ & new_n1382_ & new_n1378_ & ~new_n1376_;
  assign new_n907_ = ~new_n1401_ & ~new_n1383_ & new_n1400_ & new_n1382_ & new_n1378_ & ~new_n1376_;
  assign new_n908_ = ~new_n1401_ & ~new_n1383_ & ~new_n1400_ & ~new_n1382_ & new_n1378_ & new_n1376_;
  assign new_n909_ = ~new_n1401_ & new_n1383_ & new_n1400_ & ~new_n1382_ & new_n1378_ & new_n1376_;
  assign new_n910_ = ~new_n1401_ & ~new_n1383_ & ~new_n1400_ & new_n1382_ & new_n1378_ & new_n1376_;
  assign new_n911_ = ~new_n1401_ & new_n1383_ & ~new_n1400_ & new_n1382_ & new_n1378_ & new_n1376_;
  assign new_n912_ = ~new_n1401_ & ~new_n1383_ & new_n1400_ & new_n1382_ & new_n1378_ & new_n1376_;
  assign new_n913_ = ~new_n1401_ & new_n1383_ & new_n1400_ & new_n1382_ & new_n1378_ & new_n1376_;
  assign new_n914_ = ~new_n1401_ & new_n1383_ & ~new_n1400_ & new_n1382_ & ~new_n1378_ & ~new_n1376_;
  assign new_n915_ = new_n1401_ & ~new_n1383_ & new_n1400_ & ~new_n1382_ & new_n1378_ & ~new_n1376_;
  assign new_n916_ = new_n1401_ & ~new_n1383_ & ~new_n1400_ & new_n1382_ & new_n1378_ & ~new_n1376_;
  assign new_n917_ = new_n1401_ & new_n1383_ & ~new_n1400_ & new_n1382_ & new_n1378_ & ~new_n1376_;
  assign new_n918_ = new_n1401_ & new_n1383_ & new_n1400_ & new_n1382_ & new_n1378_ & ~new_n1376_;
  assign new_n919_ = new_n1401_ & new_n1383_ & ~new_n1400_ & ~new_n1382_ & new_n1378_ & new_n1376_;
  assign new_n920_ = ~new_n1401_ & ~new_n1383_ & ~new_n1400_ & new_n1382_ & ~new_n1378_ & ~new_n1376_;
  assign new_n921_ = new_n1401_ & new_n1383_ & new_n1400_ & ~new_n1382_ & new_n1378_ & new_n1376_;
  assign new_n922_ = new_n1401_ & ~new_n1383_ & ~new_n1400_ & new_n1382_ & new_n1378_ & new_n1376_;
  assign new_n923_ = new_n1401_ & new_n1383_ & ~new_n1400_ & new_n1382_ & new_n1378_ & new_n1376_;
  assign new_n924_ = new_n1401_ & new_n1383_ & new_n1400_ & new_n1382_ & new_n1378_ & new_n1376_;
  assign new_n925_ = ~new_n1411_ & new_n1409_ & new_n1398_ & new_n1380_ & ~new_n1397_ & new_n1381_;
  assign new_n926_ = new_n1411_ & new_n1409_ & new_n1398_ & new_n1380_ & new_n1397_ & new_n1381_;
  assign new_n927_ = new_n1411_ & ~new_n1409_ & new_n1398_ & ~new_n1380_ & ~new_n1397_ & ~new_n1381_;
  assign new_n928_ = ~new_n1396_ & ~new_n1379_ & ~new_n1427_ & ~new_n1413_ & ~new_n1377_ & ~new_n1399_;
  assign new_n929_ = ~new_n1396_ & ~new_n1379_ & new_n1427_ & ~new_n1413_ & ~new_n1377_ & ~new_n1399_;
  assign new_n930_ = new_n1401_ & new_n1383_ & new_n1400_ & ~new_n1382_ & ~new_n1378_ & ~new_n1376_;
  assign new_n931_ = ~new_n1406_ & new_n1386_ & ~new_n1404_ & ~new_n1385_ & ~new_n1384_ & ~new_n1402_;
  assign new_n932_ = ~new_n1406_ & ~new_n1386_ & new_n1404_ & ~new_n1385_ & ~new_n1384_ & ~new_n1402_;
  assign new_n933_ = ~new_n1406_ & new_n1386_ & new_n1404_ & ~new_n1385_ & ~new_n1384_ & ~new_n1402_;
  assign new_n934_ = ~new_n1406_ & new_n1386_ & ~new_n1404_ & new_n1385_ & ~new_n1384_ & ~new_n1402_;
  assign new_n935_ = ~new_n1406_ & ~new_n1386_ & new_n1404_ & new_n1385_ & ~new_n1384_ & ~new_n1402_;
  assign new_n936_ = ~new_n1406_ & new_n1386_ & new_n1404_ & new_n1385_ & ~new_n1384_ & ~new_n1402_;
  assign new_n937_ = ~new_n1406_ & new_n1386_ & new_n1404_ & ~new_n1385_ & ~new_n1384_ & new_n1402_;
  assign new_n938_ = ~new_n1406_ & ~new_n1386_ & ~new_n1404_ & new_n1385_ & ~new_n1384_ & new_n1402_;
  assign new_n939_ = ~new_n1406_ & new_n1386_ & ~new_n1404_ & new_n1385_ & ~new_n1384_ & new_n1402_;
  assign new_n940_ = ~new_n1406_ & new_n1386_ & new_n1404_ & new_n1385_ & ~new_n1384_ & new_n1402_;
  assign new_n941_ = new_n1406_ & ~new_n1386_ & ~new_n1404_ & ~new_n1385_ & ~new_n1384_ & ~new_n1402_;
  assign new_n942_ = new_n1406_ & ~new_n1386_ & new_n1404_ & ~new_n1385_ & ~new_n1384_ & ~new_n1402_;
  assign new_n943_ = new_n1406_ & new_n1386_ & new_n1404_ & ~new_n1385_ & ~new_n1384_ & ~new_n1402_;
  assign new_n944_ = new_n1406_ & ~new_n1386_ & ~new_n1404_ & new_n1385_ & ~new_n1384_ & ~new_n1402_;
  assign new_n945_ = new_n1406_ & new_n1386_ & ~new_n1404_ & new_n1385_ & ~new_n1384_ & ~new_n1402_;
  assign new_n946_ = new_n1406_ & new_n1386_ & new_n1404_ & new_n1385_ & ~new_n1384_ & ~new_n1402_;
  assign new_n947_ = new_n1406_ & new_n1386_ & ~new_n1404_ & ~new_n1385_ & ~new_n1384_ & new_n1402_;
  assign new_n948_ = new_n1406_ & new_n1386_ & new_n1404_ & ~new_n1385_ & ~new_n1384_ & new_n1402_;
  assign new_n949_ = new_n1406_ & ~new_n1386_ & new_n1404_ & new_n1385_ & ~new_n1384_ & new_n1402_;
  assign new_n950_ = new_n1406_ & new_n1386_ & new_n1404_ & new_n1385_ & ~new_n1384_ & new_n1402_;
  assign new_n951_ = ~new_n1406_ & ~new_n1386_ & ~new_n1404_ & ~new_n1385_ & new_n1384_ & ~new_n1402_;
  assign new_n952_ = ~new_n1406_ & new_n1386_ & ~new_n1404_ & ~new_n1385_ & new_n1384_ & ~new_n1402_;
  assign new_n953_ = ~new_n1406_ & ~new_n1386_ & new_n1404_ & ~new_n1385_ & new_n1384_ & ~new_n1402_;
  assign new_n954_ = ~new_n1406_ & ~new_n1386_ & ~new_n1404_ & new_n1385_ & new_n1384_ & ~new_n1402_;
  assign new_n955_ = ~new_n1406_ & new_n1386_ & ~new_n1404_ & new_n1385_ & new_n1384_ & ~new_n1402_;
  assign new_n956_ = ~new_n1406_ & ~new_n1386_ & new_n1404_ & new_n1385_ & new_n1384_ & ~new_n1402_;
  assign new_n957_ = ~new_n1406_ & new_n1386_ & new_n1404_ & new_n1385_ & new_n1384_ & ~new_n1402_;
  assign new_n958_ = ~new_n1406_ & ~new_n1386_ & ~new_n1404_ & ~new_n1385_ & new_n1384_ & new_n1402_;
  assign new_n959_ = ~new_n1406_ & ~new_n1386_ & new_n1404_ & ~new_n1385_ & new_n1384_ & new_n1402_;
  assign new_n960_ = ~new_n1406_ & new_n1386_ & new_n1404_ & ~new_n1385_ & new_n1384_ & new_n1402_;
  assign new_n961_ = ~new_n1406_ & ~new_n1386_ & ~new_n1404_ & new_n1385_ & new_n1384_ & new_n1402_;
  assign new_n962_ = new_n1406_ & ~new_n1386_ & ~new_n1404_ & ~new_n1385_ & new_n1384_ & ~new_n1402_;
  assign new_n963_ = new_n1406_ & new_n1386_ & ~new_n1404_ & ~new_n1385_ & new_n1384_ & ~new_n1402_;
  assign new_n964_ = new_n1406_ & new_n1386_ & new_n1404_ & ~new_n1385_ & new_n1384_ & ~new_n1402_;
  assign new_n965_ = new_n1406_ & ~new_n1386_ & ~new_n1404_ & new_n1385_ & new_n1384_ & ~new_n1402_;
  assign new_n966_ = new_n1406_ & ~new_n1386_ & new_n1404_ & new_n1385_ & new_n1384_ & ~new_n1402_;
  assign new_n967_ = new_n1406_ & ~new_n1386_ & ~new_n1404_ & ~new_n1385_ & new_n1384_ & new_n1402_;
  assign new_n968_ = new_n1406_ & ~new_n1386_ & new_n1404_ & ~new_n1385_ & new_n1384_ & new_n1402_;
  assign new_n969_ = new_n1406_ & new_n1386_ & new_n1404_ & ~new_n1385_ & new_n1384_ & new_n1402_;
  assign new_n970_ = new_n1406_ & ~new_n1386_ & ~new_n1404_ & new_n1385_ & new_n1384_ & new_n1402_;
  assign new_n971_ = new_n1406_ & new_n1386_ & ~new_n1404_ & new_n1385_ & new_n1384_ & new_n1402_;
  assign new_n972_ = new_n1406_ & new_n1386_ & new_n1404_ & new_n1385_ & new_n1384_ & new_n1402_;
  assign new_n973_ = ~new_n1411_ & new_n1409_ & ~new_n1398_ & new_n1380_ & ~new_n1397_ & new_n1381_;
  assign new_n974_ = new_n1396_ & new_n1379_ & ~new_n1427_ & ~new_n1413_ & ~new_n1377_ & ~new_n1399_;
  assign new_n975_ = ~new_n1396_ & new_n1379_ & ~new_n1427_ & ~new_n1413_ & new_n1377_ & ~new_n1399_;
  assign new_n976_ = new_n1401_ & new_n1383_ & ~new_n1400_ & ~new_n1382_ & new_n1378_ & ~new_n1376_;
  assign new_n977_ = ~new_n1390_ & new_n1389_ & ~new_n1410_ & ~new_n1388_ & ~new_n1387_ & ~new_n1408_;
  assign new_n978_ = ~new_n1390_ & ~new_n1389_ & ~new_n1410_ & new_n1388_ & ~new_n1387_ & ~new_n1408_;
  assign new_n979_ = ~new_n1390_ & new_n1389_ & ~new_n1410_ & new_n1388_ & ~new_n1387_ & ~new_n1408_;
  assign new_n980_ = ~new_n1390_ & ~new_n1389_ & new_n1410_ & new_n1388_ & ~new_n1387_ & ~new_n1408_;
  assign new_n981_ = ~new_n1390_ & new_n1389_ & new_n1410_ & new_n1388_ & ~new_n1387_ & ~new_n1408_;
  assign new_n982_ = ~new_n1390_ & new_n1389_ & ~new_n1410_ & ~new_n1388_ & ~new_n1387_ & new_n1408_;
  assign new_n983_ = ~new_n1390_ & ~new_n1389_ & new_n1410_ & ~new_n1388_ & ~new_n1387_ & new_n1408_;
  assign new_n984_ = ~new_n1390_ & new_n1389_ & new_n1410_ & ~new_n1388_ & ~new_n1387_ & new_n1408_;
  assign new_n985_ = ~new_n1390_ & ~new_n1389_ & ~new_n1410_ & new_n1388_ & ~new_n1387_ & new_n1408_;
  assign new_n986_ = ~new_n1390_ & ~new_n1389_ & new_n1410_ & new_n1388_ & ~new_n1387_ & new_n1408_;
  assign new_n987_ = ~new_n1390_ & new_n1389_ & new_n1410_ & new_n1388_ & ~new_n1387_ & new_n1408_;
  assign new_n988_ = new_n1390_ & ~new_n1389_ & ~new_n1410_ & ~new_n1388_ & ~new_n1387_ & ~new_n1408_;
  assign new_n989_ = new_n1390_ & new_n1389_ & ~new_n1410_ & ~new_n1388_ & ~new_n1387_ & ~new_n1408_;
  assign new_n990_ = new_n1390_ & new_n1389_ & new_n1410_ & ~new_n1388_ & ~new_n1387_ & ~new_n1408_;
  assign new_n991_ = new_n1390_ & new_n1389_ & ~new_n1410_ & new_n1388_ & ~new_n1387_ & ~new_n1408_;
  assign new_n992_ = new_n1390_ & ~new_n1389_ & new_n1410_ & new_n1388_ & ~new_n1387_ & ~new_n1408_;
  assign new_n993_ = new_n1390_ & ~new_n1389_ & ~new_n1410_ & ~new_n1388_ & ~new_n1387_ & new_n1408_;
  assign new_n994_ = new_n1401_ & ~new_n1383_ & new_n1400_ & ~new_n1382_ & new_n1378_ & new_n1376_;
  assign new_n995_ = new_n1390_ & new_n1389_ & new_n1410_ & ~new_n1388_ & ~new_n1387_ & new_n1408_;
  assign new_n996_ = new_n1390_ & ~new_n1389_ & ~new_n1410_ & new_n1388_ & ~new_n1387_ & new_n1408_;
  assign new_n997_ = new_n1390_ & new_n1389_ & ~new_n1410_ & new_n1388_ & ~new_n1387_ & new_n1408_;
  assign new_n998_ = new_n1390_ & new_n1389_ & new_n1410_ & new_n1388_ & ~new_n1387_ & new_n1408_;
  assign new_n999_ = ~new_n1390_ & new_n1389_ & new_n1410_ & ~new_n1388_ & new_n1387_ & ~new_n1408_;
  assign new_n1000_ = ~new_n1390_ & ~new_n1389_ & ~new_n1410_ & new_n1388_ & new_n1387_ & ~new_n1408_;
  assign new_n1001_ = ~new_n1390_ & new_n1389_ & ~new_n1410_ & new_n1388_ & new_n1387_ & ~new_n1408_;
  assign new_n1002_ = ~new_n1390_ & ~new_n1389_ & new_n1410_ & new_n1388_ & new_n1387_ & ~new_n1408_;
  assign new_n1003_ = ~new_n1390_ & ~new_n1389_ & ~new_n1410_ & ~new_n1388_ & new_n1387_ & new_n1408_;
  assign new_n1004_ = ~new_n1390_ & new_n1389_ & ~new_n1410_ & ~new_n1388_ & new_n1387_ & new_n1408_;
  assign new_n1005_ = ~new_n1411_ & ~new_n1409_ & ~new_n1398_ & new_n1380_ & ~new_n1397_ & new_n1381_;
  assign new_n1006_ = ~new_n1390_ & ~new_n1389_ & ~new_n1410_ & new_n1388_ & new_n1387_ & new_n1408_;
  assign new_n1007_ = ~new_n1390_ & new_n1389_ & ~new_n1410_ & new_n1388_ & new_n1387_ & new_n1408_;
  assign new_n1008_ = ~new_n1390_ & new_n1389_ & new_n1410_ & new_n1388_ & new_n1387_ & new_n1408_;
  assign new_n1009_ = new_n1390_ & ~new_n1389_ & ~new_n1410_ & ~new_n1388_ & new_n1387_ & ~new_n1408_;
  assign new_n1010_ = new_n1390_ & ~new_n1389_ & new_n1410_ & ~new_n1388_ & new_n1387_ & ~new_n1408_;
  assign new_n1011_ = new_n1390_ & new_n1389_ & new_n1410_ & ~new_n1388_ & new_n1387_ & ~new_n1408_;
  assign new_n1012_ = new_n1390_ & new_n1389_ & ~new_n1410_ & new_n1388_ & new_n1387_ & ~new_n1408_;
  assign new_n1013_ = new_n1390_ & new_n1389_ & new_n1410_ & new_n1388_ & new_n1387_ & ~new_n1408_;
  assign new_n1014_ = new_n1390_ & ~new_n1389_ & ~new_n1410_ & ~new_n1388_ & new_n1387_ & new_n1408_;
  assign new_n1015_ = new_n1390_ & new_n1389_ & ~new_n1410_ & ~new_n1388_ & new_n1387_ & new_n1408_;
  assign new_n1016_ = new_n1390_ & new_n1389_ & new_n1410_ & ~new_n1388_ & new_n1387_ & new_n1408_;
  assign new_n1017_ = new_n1390_ & ~new_n1389_ & ~new_n1410_ & new_n1388_ & new_n1387_ & new_n1408_;
  assign new_n1018_ = new_n1390_ & ~new_n1389_ & new_n1410_ & new_n1388_ & new_n1387_ & new_n1408_;
  assign new_n1019_ = new_n1390_ & new_n1389_ & new_n1410_ & new_n1388_ & new_n1387_ & new_n1408_;
  assign new_n1020_ = ~new_n1411_ & new_n1409_ & new_n1398_ & ~new_n1380_ & ~new_n1397_ & new_n1381_;
  assign new_n1021_ = ~new_n1396_ & new_n1379_ & ~new_n1427_ & ~new_n1413_ & ~new_n1377_ & ~new_n1399_;
  assign new_n1022_ = new_n1396_ & ~new_n1379_ & ~new_n1427_ & ~new_n1413_ & new_n1377_ & ~new_n1399_;
  assign new_n1023_ = ~new_n1406_ & ~new_n1386_ & ~new_n1404_ & ~new_n1385_ & ~new_n1384_ & ~new_n1402_;
  assign new_n1024_ = ~new_n1394_ & ~new_n1393_ & ~new_n1414_ & ~new_n1392_ & ~new_n1412_ & ~new_n1391_;
  assign new_n1025_ = ~new_n1394_ & ~new_n1393_ & new_n1414_ & ~new_n1392_ & ~new_n1412_ & ~new_n1391_;
  assign new_n1026_ = ~new_n1394_ & new_n1393_ & new_n1414_ & ~new_n1392_ & ~new_n1412_ & ~new_n1391_;
  assign new_n1027_ = ~new_n1394_ & ~new_n1393_ & ~new_n1414_ & new_n1392_ & ~new_n1412_ & ~new_n1391_;
  assign new_n1028_ = ~new_n1394_ & ~new_n1393_ & new_n1414_ & new_n1392_ & ~new_n1412_ & ~new_n1391_;
  assign new_n1029_ = new_n1406_ & new_n1386_ & ~new_n1404_ & new_n1385_ & ~new_n1384_ & new_n1402_;
  assign new_n1030_ = ~new_n1394_ & ~new_n1393_ & new_n1414_ & ~new_n1392_ & ~new_n1412_ & new_n1391_;
  assign new_n1031_ = ~new_n1394_ & ~new_n1393_ & ~new_n1414_ & new_n1392_ & ~new_n1412_ & new_n1391_;
  assign new_n1032_ = ~new_n1394_ & new_n1393_ & ~new_n1414_ & new_n1392_ & ~new_n1412_ & new_n1391_;
  assign new_n1033_ = ~new_n1394_ & ~new_n1393_ & new_n1414_ & new_n1392_ & ~new_n1412_ & new_n1391_;
  assign new_n1034_ = ~new_n1394_ & new_n1393_ & new_n1414_ & new_n1392_ & ~new_n1412_ & new_n1391_;
  assign new_n1035_ = new_n1394_ & ~new_n1393_ & ~new_n1414_ & ~new_n1392_ & ~new_n1412_ & ~new_n1391_;
  assign new_n1036_ = new_n1394_ & new_n1393_ & ~new_n1414_ & ~new_n1392_ & ~new_n1412_ & ~new_n1391_;
  assign new_n1037_ = new_n1394_ & ~new_n1393_ & ~new_n1414_ & new_n1392_ & ~new_n1412_ & ~new_n1391_;
  assign new_n1038_ = new_n1394_ & new_n1393_ & ~new_n1414_ & new_n1392_ & ~new_n1412_ & ~new_n1391_;
  assign new_n1039_ = new_n1394_ & ~new_n1393_ & new_n1414_ & new_n1392_ & ~new_n1412_ & ~new_n1391_;
  assign new_n1040_ = new_n1394_ & new_n1393_ & new_n1414_ & new_n1392_ & ~new_n1412_ & ~new_n1391_;
  assign new_n1041_ = new_n1394_ & ~new_n1393_ & ~new_n1414_ & ~new_n1392_ & ~new_n1412_ & new_n1391_;
  assign new_n1042_ = new_n1394_ & ~new_n1393_ & new_n1414_ & ~new_n1392_ & ~new_n1412_ & new_n1391_;
  assign new_n1043_ = new_n1394_ & new_n1393_ & new_n1414_ & ~new_n1392_ & ~new_n1412_ & new_n1391_;
  assign new_n1044_ = new_n1394_ & new_n1393_ & ~new_n1414_ & new_n1392_ & ~new_n1412_ & new_n1391_;
  assign new_n1045_ = new_n1394_ & ~new_n1393_ & new_n1414_ & new_n1392_ & ~new_n1412_ & new_n1391_;
  assign new_n1046_ = ~new_n1394_ & ~new_n1393_ & ~new_n1414_ & ~new_n1392_ & new_n1412_ & ~new_n1391_;
  assign new_n1047_ = ~new_n1394_ & new_n1393_ & ~new_n1414_ & ~new_n1392_ & new_n1412_ & ~new_n1391_;
  assign new_n1048_ = ~new_n1394_ & ~new_n1393_ & new_n1414_ & ~new_n1392_ & new_n1412_ & ~new_n1391_;
  assign new_n1049_ = ~new_n1394_ & new_n1393_ & new_n1414_ & ~new_n1392_ & new_n1412_ & ~new_n1391_;
  assign new_n1050_ = ~new_n1394_ & ~new_n1393_ & new_n1414_ & new_n1392_ & new_n1412_ & ~new_n1391_;
  assign new_n1051_ = ~new_n1394_ & new_n1393_ & new_n1414_ & new_n1392_ & new_n1412_ & ~new_n1391_;
  assign new_n1052_ = ~new_n1394_ & ~new_n1393_ & ~new_n1414_ & ~new_n1392_ & new_n1412_ & new_n1391_;
  assign new_n1053_ = ~new_n1394_ & new_n1393_ & new_n1414_ & ~new_n1392_ & new_n1412_ & new_n1391_;
  assign new_n1054_ = ~new_n1394_ & new_n1393_ & ~new_n1414_ & new_n1392_ & new_n1412_ & new_n1391_;
  assign new_n1055_ = ~new_n1394_ & ~new_n1393_ & new_n1414_ & new_n1392_ & new_n1412_ & new_n1391_;
  assign new_n1056_ = ~new_n1394_ & new_n1393_ & new_n1414_ & new_n1392_ & new_n1412_ & new_n1391_;
  assign new_n1057_ = new_n1394_ & new_n1393_ & ~new_n1414_ & ~new_n1392_ & new_n1412_ & ~new_n1391_;
  assign new_n1058_ = new_n1394_ & new_n1393_ & new_n1414_ & ~new_n1392_ & new_n1412_ & ~new_n1391_;
  assign new_n1059_ = new_n1394_ & ~new_n1393_ & ~new_n1414_ & new_n1392_ & new_n1412_ & ~new_n1391_;
  assign new_n1060_ = new_n1394_ & new_n1393_ & ~new_n1414_ & new_n1392_ & new_n1412_ & ~new_n1391_;
  assign new_n1061_ = new_n1394_ & ~new_n1393_ & new_n1414_ & new_n1392_ & new_n1412_ & ~new_n1391_;
  assign new_n1062_ = new_n1394_ & new_n1393_ & new_n1414_ & new_n1392_ & new_n1412_ & ~new_n1391_;
  assign new_n1063_ = new_n1394_ & ~new_n1393_ & ~new_n1414_ & ~new_n1392_ & new_n1412_ & new_n1391_;
  assign new_n1064_ = new_n1394_ & new_n1393_ & ~new_n1414_ & ~new_n1392_ & new_n1412_ & new_n1391_;
  assign new_n1065_ = ~new_n1411_ & ~new_n1409_ & new_n1398_ & ~new_n1380_ & ~new_n1397_ & new_n1381_;
  assign new_n1066_ = new_n1394_ & new_n1393_ & new_n1414_ & ~new_n1392_ & new_n1412_ & new_n1391_;
  assign new_n1067_ = new_n1394_ & ~new_n1393_ & ~new_n1414_ & new_n1392_ & new_n1412_ & new_n1391_;
  assign new_n1068_ = new_n1394_ & new_n1393_ & new_n1414_ & new_n1392_ & new_n1412_ & new_n1391_;
  assign new_n1069_ = ~new_n1411_ & new_n1409_ & ~new_n1398_ & ~new_n1380_ & ~new_n1397_ & new_n1381_;
  assign new_n1070_ = new_n1411_ & ~new_n1409_ & new_n1398_ & new_n1380_ & new_n1397_ & new_n1381_;
  assign new_n1071_ = new_n1411_ & ~new_n1409_ & ~new_n1398_ & new_n1380_ & new_n1397_ & new_n1381_;
  assign new_n1072_ = new_n1411_ & new_n1409_ & new_n1398_ & ~new_n1380_ & new_n1397_ & new_n1381_;
  assign new_n1073_ = ~new_n1420_ & new_n1419_ & ~new_n1418_ & ~new_n1417_ & ~new_n1415_ & ~new_n1416_;
  assign new_n1074_ = ~new_n1420_ & new_n1419_ & new_n1418_ & ~new_n1417_ & ~new_n1415_ & ~new_n1416_;
  assign new_n1075_ = ~new_n1420_ & ~new_n1419_ & ~new_n1418_ & new_n1417_ & ~new_n1415_ & ~new_n1416_;
  assign new_n1076_ = ~new_n1420_ & new_n1419_ & new_n1418_ & new_n1417_ & ~new_n1415_ & ~new_n1416_;
  assign new_n1077_ = ~new_n1420_ & ~new_n1419_ & ~new_n1418_ & ~new_n1417_ & ~new_n1415_ & new_n1416_;
  assign new_n1078_ = ~new_n1420_ & new_n1419_ & ~new_n1418_ & ~new_n1417_ & ~new_n1415_ & new_n1416_;
  assign new_n1079_ = ~new_n1420_ & ~new_n1419_ & new_n1418_ & ~new_n1417_ & ~new_n1415_ & new_n1416_;
  assign new_n1080_ = ~new_n1420_ & new_n1419_ & new_n1418_ & ~new_n1417_ & ~new_n1415_ & new_n1416_;
  assign new_n1081_ = ~new_n1420_ & ~new_n1419_ & ~new_n1418_ & new_n1417_ & ~new_n1415_ & new_n1416_;
  assign new_n1082_ = ~new_n1420_ & new_n1419_ & ~new_n1418_ & new_n1417_ & ~new_n1415_ & new_n1416_;
  assign new_n1083_ = ~new_n1420_ & ~new_n1419_ & new_n1418_ & new_n1417_ & ~new_n1415_ & new_n1416_;
  assign new_n1084_ = new_n1420_ & ~new_n1419_ & ~new_n1418_ & ~new_n1417_ & ~new_n1415_ & ~new_n1416_;
  assign new_n1085_ = new_n1420_ & ~new_n1419_ & new_n1418_ & ~new_n1417_ & ~new_n1415_ & ~new_n1416_;
  assign new_n1086_ = new_n1420_ & new_n1419_ & new_n1418_ & ~new_n1417_ & ~new_n1415_ & ~new_n1416_;
  assign new_n1087_ = new_n1420_ & new_n1419_ & ~new_n1418_ & new_n1417_ & ~new_n1415_ & ~new_n1416_;
  assign new_n1088_ = new_n1420_ & new_n1419_ & new_n1418_ & new_n1417_ & ~new_n1415_ & ~new_n1416_;
  assign new_n1089_ = new_n1420_ & ~new_n1419_ & ~new_n1418_ & ~new_n1417_ & ~new_n1415_ & new_n1416_;
  assign new_n1090_ = new_n1420_ & new_n1419_ & ~new_n1418_ & ~new_n1417_ & ~new_n1415_ & new_n1416_;
  assign new_n1091_ = new_n1420_ & ~new_n1419_ & new_n1418_ & ~new_n1417_ & ~new_n1415_ & new_n1416_;
  assign new_n1092_ = new_n1420_ & new_n1419_ & new_n1418_ & ~new_n1417_ & ~new_n1415_ & new_n1416_;
  assign new_n1093_ = new_n1420_ & new_n1419_ & ~new_n1418_ & new_n1417_ & ~new_n1415_ & new_n1416_;
  assign new_n1094_ = new_n1420_ & new_n1419_ & new_n1418_ & new_n1417_ & ~new_n1415_ & new_n1416_;
  assign new_n1095_ = ~new_n1420_ & ~new_n1419_ & new_n1418_ & ~new_n1417_ & new_n1415_ & ~new_n1416_;
  assign new_n1096_ = ~new_n1420_ & new_n1419_ & new_n1418_ & ~new_n1417_ & new_n1415_ & ~new_n1416_;
  assign new_n1097_ = ~new_n1420_ & ~new_n1419_ & ~new_n1418_ & new_n1417_ & new_n1415_ & ~new_n1416_;
  assign new_n1098_ = ~new_n1420_ & new_n1419_ & ~new_n1418_ & new_n1417_ & new_n1415_ & ~new_n1416_;
  assign new_n1099_ = ~new_n1420_ & ~new_n1419_ & new_n1418_ & new_n1417_ & new_n1415_ & ~new_n1416_;
  assign new_n1100_ = ~new_n1420_ & new_n1419_ & new_n1418_ & new_n1417_ & new_n1415_ & ~new_n1416_;
  assign new_n1101_ = ~new_n1420_ & ~new_n1419_ & ~new_n1418_ & ~new_n1417_ & new_n1415_ & new_n1416_;
  assign new_n1102_ = ~new_n1420_ & new_n1419_ & ~new_n1418_ & ~new_n1417_ & new_n1415_ & new_n1416_;
  assign new_n1103_ = ~new_n1420_ & ~new_n1419_ & new_n1418_ & ~new_n1417_ & new_n1415_ & new_n1416_;
  assign new_n1104_ = ~new_n1420_ & new_n1419_ & ~new_n1418_ & new_n1417_ & new_n1415_ & new_n1416_;
  assign new_n1105_ = ~new_n1420_ & ~new_n1419_ & new_n1418_ & new_n1417_ & new_n1415_ & new_n1416_;
  assign new_n1106_ = new_n1420_ & ~new_n1419_ & ~new_n1418_ & ~new_n1417_ & new_n1415_ & ~new_n1416_;
  assign new_n1107_ = new_n1420_ & new_n1419_ & ~new_n1418_ & ~new_n1417_ & new_n1415_ & ~new_n1416_;
  assign new_n1108_ = new_n1420_ & ~new_n1419_ & new_n1418_ & ~new_n1417_ & new_n1415_ & ~new_n1416_;
  assign new_n1109_ = new_n1420_ & ~new_n1419_ & new_n1418_ & new_n1417_ & new_n1415_ & ~new_n1416_;
  assign new_n1110_ = new_n1420_ & new_n1419_ & new_n1418_ & new_n1417_ & new_n1415_ & ~new_n1416_;
  assign new_n1111_ = new_n1420_ & ~new_n1419_ & ~new_n1418_ & ~new_n1417_ & new_n1415_ & new_n1416_;
  assign new_n1112_ = new_n1420_ & new_n1419_ & ~new_n1418_ & ~new_n1417_ & new_n1415_ & new_n1416_;
  assign new_n1113_ = new_n1420_ & new_n1419_ & new_n1418_ & ~new_n1417_ & new_n1415_ & new_n1416_;
  assign new_n1114_ = new_n1420_ & ~new_n1419_ & ~new_n1418_ & new_n1417_ & new_n1415_ & new_n1416_;
  assign new_n1115_ = new_n1420_ & ~new_n1419_ & new_n1418_ & new_n1417_ & new_n1415_ & new_n1416_;
  assign new_n1116_ = new_n1420_ & new_n1419_ & new_n1418_ & new_n1417_ & new_n1415_ & new_n1416_;
  assign new_n1117_ = ~new_n1411_ & ~new_n1409_ & ~new_n1398_ & ~new_n1380_ & ~new_n1397_ & new_n1381_;
  assign new_n1118_ = new_n1411_ & ~new_n1409_ & new_n1398_ & ~new_n1380_ & new_n1397_ & new_n1381_;
  assign new_n1119_ = new_n1411_ & new_n1409_ & ~new_n1398_ & ~new_n1380_ & new_n1397_ & new_n1381_;
  assign new_n1120_ = new_n1411_ & ~new_n1409_ & ~new_n1398_ & ~new_n1380_ & new_n1397_ & new_n1381_;
  assign new_n1121_ = ~new_n1426_ & ~new_n1425_ & ~new_n1424_ & ~new_n1423_ & ~new_n1421_ & ~new_n1422_;
  assign new_n1122_ = ~new_n1426_ & ~new_n1425_ & ~new_n1424_ & new_n1423_ & ~new_n1421_ & ~new_n1422_;
  assign new_n1123_ = ~new_n1426_ & new_n1425_ & ~new_n1424_ & new_n1423_ & ~new_n1421_ & ~new_n1422_;
  assign new_n1124_ = ~new_n1426_ & ~new_n1425_ & new_n1424_ & new_n1423_ & ~new_n1421_ & ~new_n1422_;
  assign new_n1125_ = ~new_n1426_ & ~new_n1425_ & ~new_n1424_ & ~new_n1423_ & ~new_n1421_ & new_n1422_;
  assign new_n1126_ = ~new_n1426_ & new_n1425_ & ~new_n1424_ & ~new_n1423_ & ~new_n1421_ & new_n1422_;
  assign new_n1127_ = ~new_n1426_ & ~new_n1425_ & new_n1424_ & ~new_n1423_ & ~new_n1421_ & new_n1422_;
  assign new_n1128_ = ~new_n1426_ & new_n1425_ & new_n1424_ & ~new_n1423_ & ~new_n1421_ & new_n1422_;
  assign new_n1129_ = ~new_n1426_ & ~new_n1425_ & ~new_n1424_ & new_n1423_ & ~new_n1421_ & new_n1422_;
  assign new_n1130_ = ~new_n1426_ & ~new_n1425_ & new_n1424_ & new_n1423_ & ~new_n1421_ & new_n1422_;
  assign new_n1131_ = ~new_n1426_ & new_n1425_ & new_n1424_ & new_n1423_ & ~new_n1421_ & new_n1422_;
  assign new_n1132_ = new_n1426_ & new_n1425_ & ~new_n1424_ & ~new_n1423_ & ~new_n1421_ & ~new_n1422_;
  assign new_n1133_ = new_n1426_ & ~new_n1425_ & new_n1424_ & ~new_n1423_ & ~new_n1421_ & ~new_n1422_;
  assign new_n1134_ = new_n1426_ & ~new_n1425_ & ~new_n1424_ & new_n1423_ & ~new_n1421_ & ~new_n1422_;
  assign new_n1135_ = new_n1426_ & new_n1425_ & ~new_n1424_ & new_n1423_ & ~new_n1421_ & ~new_n1422_;
  assign new_n1136_ = new_n1426_ & ~new_n1425_ & new_n1424_ & new_n1423_ & ~new_n1421_ & ~new_n1422_;
  assign new_n1137_ = new_n1426_ & ~new_n1425_ & ~new_n1424_ & ~new_n1423_ & ~new_n1421_ & new_n1422_;
  assign new_n1138_ = new_n1426_ & new_n1425_ & ~new_n1424_ & ~new_n1423_ & ~new_n1421_ & new_n1422_;
  assign new_n1139_ = new_n1426_ & ~new_n1425_ & new_n1424_ & ~new_n1423_ & ~new_n1421_ & new_n1422_;
  assign new_n1140_ = new_n1426_ & new_n1425_ & new_n1424_ & ~new_n1423_ & ~new_n1421_ & new_n1422_;
  assign new_n1141_ = new_n1426_ & new_n1425_ & ~new_n1424_ & new_n1423_ & ~new_n1421_ & new_n1422_;
  assign new_n1142_ = new_n1426_ & ~new_n1425_ & new_n1424_ & new_n1423_ & ~new_n1421_ & new_n1422_;
  assign new_n1143_ = ~new_n1426_ & ~new_n1425_ & ~new_n1424_ & ~new_n1423_ & new_n1421_ & ~new_n1422_;
  assign new_n1144_ = ~new_n1426_ & new_n1425_ & ~new_n1424_ & ~new_n1423_ & new_n1421_ & ~new_n1422_;
  assign new_n1145_ = ~new_n1426_ & ~new_n1425_ & ~new_n1424_ & new_n1423_ & new_n1421_ & ~new_n1422_;
  assign new_n1146_ = ~new_n1426_ & new_n1425_ & ~new_n1424_ & new_n1423_ & new_n1421_ & ~new_n1422_;
  assign new_n1147_ = ~new_n1426_ & ~new_n1425_ & new_n1424_ & new_n1423_ & new_n1421_ & ~new_n1422_;
  assign new_n1148_ = ~new_n1426_ & new_n1425_ & ~new_n1424_ & ~new_n1423_ & new_n1421_ & new_n1422_;
  assign new_n1149_ = ~new_n1426_ & ~new_n1425_ & new_n1424_ & ~new_n1423_ & new_n1421_ & new_n1422_;
  assign new_n1150_ = ~new_n1426_ & new_n1425_ & new_n1424_ & ~new_n1423_ & new_n1421_ & new_n1422_;
  assign new_n1151_ = ~new_n1426_ & ~new_n1425_ & ~new_n1424_ & new_n1423_ & new_n1421_ & new_n1422_;
  assign new_n1152_ = ~new_n1426_ & new_n1425_ & ~new_n1424_ & new_n1423_ & new_n1421_ & new_n1422_;
  assign new_n1153_ = ~new_n1426_ & ~new_n1425_ & new_n1424_ & new_n1423_ & new_n1421_ & new_n1422_;
  assign new_n1154_ = new_n1426_ & ~new_n1425_ & new_n1424_ & ~new_n1423_ & new_n1421_ & ~new_n1422_;
  assign new_n1155_ = new_n1426_ & new_n1425_ & new_n1424_ & ~new_n1423_ & new_n1421_ & ~new_n1422_;
  assign new_n1156_ = new_n1426_ & new_n1425_ & ~new_n1424_ & new_n1423_ & new_n1421_ & ~new_n1422_;
  assign new_n1157_ = new_n1426_ & new_n1425_ & new_n1424_ & new_n1423_ & new_n1421_ & ~new_n1422_;
  assign new_n1158_ = new_n1426_ & ~new_n1425_ & ~new_n1424_ & ~new_n1423_ & new_n1421_ & new_n1422_;
  assign new_n1159_ = new_n1426_ & new_n1425_ & ~new_n1424_ & ~new_n1423_ & new_n1421_ & new_n1422_;
  assign new_n1160_ = new_n1426_ & ~new_n1425_ & new_n1424_ & ~new_n1423_ & new_n1421_ & new_n1422_;
  assign new_n1161_ = new_n1426_ & ~new_n1425_ & ~new_n1424_ & new_n1423_ & new_n1421_ & new_n1422_;
  assign new_n1162_ = new_n1426_ & new_n1425_ & ~new_n1424_ & new_n1423_ & new_n1421_ & new_n1422_;
  assign new_n1163_ = new_n1426_ & ~new_n1425_ & new_n1424_ & new_n1423_ & new_n1421_ & new_n1422_;
  assign new_n1164_ = new_n1426_ & new_n1425_ & new_n1424_ & new_n1423_ & new_n1421_ & new_n1422_;
  assign new_n1165_ = new_n1411_ & new_n1409_ & new_n1398_ & new_n1380_ & new_n1397_ & ~new_n1381_;
  assign new_n1166_ = new_n1411_ & new_n1409_ & ~new_n1398_ & new_n1380_ & new_n1397_ & ~new_n1381_;
  assign new_n1167_ = ~new_n1390_ & ~new_n1389_ & new_n1410_ & ~new_n1388_ & new_n1387_ & new_n1408_;
  assign new_n1168_ = new_n1411_ & new_n1409_ & ~new_n1398_ & ~new_n1380_ & new_n1397_ & ~new_n1381_;
  assign new_n1169_ = new_n1411_ & ~new_n1409_ & ~new_n1398_ & ~new_n1380_ & new_n1397_ & ~new_n1381_;
  assign new_n1170_ = ~new_n1411_ & ~new_n1409_ & new_n1398_ & new_n1380_ & new_n1397_ & new_n1381_;
  assign new_n1171_ = ~new_n1411_ & new_n1409_ & ~new_n1398_ & new_n1380_ & new_n1397_ & new_n1381_;
  assign new_n1172_ = ~new_n1411_ & ~new_n1409_ & ~new_n1398_ & new_n1380_ & new_n1397_ & new_n1381_;
  assign new_n1173_ = ~new_n1411_ & new_n1409_ & new_n1398_ & ~new_n1380_ & new_n1397_ & new_n1381_;
  assign new_n1174_ = ~new_n1411_ & ~new_n1409_ & new_n1398_ & ~new_n1380_ & new_n1397_ & new_n1381_;
  assign new_n1175_ = ~new_n1411_ & new_n1409_ & ~new_n1398_ & ~new_n1380_ & new_n1397_ & new_n1381_;
  assign new_n1176_ = ~new_n1411_ & ~new_n1409_ & ~new_n1398_ & ~new_n1380_ & new_n1397_ & new_n1381_;
  assign new_n1177_ = ~new_n1411_ & new_n1409_ & new_n1398_ & new_n1380_ & new_n1397_ & ~new_n1381_;
  assign new_n1178_ = ~new_n1411_ & new_n1409_ & ~new_n1398_ & new_n1380_ & new_n1397_ & ~new_n1381_;
  assign new_n1179_ = ~new_n1411_ & ~new_n1409_ & ~new_n1398_ & new_n1380_ & new_n1397_ & ~new_n1381_;
  assign new_n1180_ = ~new_n1411_ & ~new_n1409_ & new_n1398_ & ~new_n1380_ & new_n1397_ & ~new_n1381_;
  assign new_n1181_ = new_n1411_ & ~new_n1409_ & new_n1398_ & new_n1380_ & ~new_n1397_ & new_n1381_;
  assign new_n1182_ = new_n1411_ & new_n1409_ & ~new_n1398_ & new_n1380_ & ~new_n1397_ & new_n1381_;
  assign new_n1183_ = new_n1411_ & ~new_n1409_ & ~new_n1398_ & new_n1380_ & ~new_n1397_ & new_n1381_;
  assign new_n1184_ = new_n1411_ & new_n1409_ & new_n1398_ & ~new_n1380_ & ~new_n1397_ & new_n1381_;
  assign new_n1185_ = new_n1411_ & ~new_n1409_ & new_n1398_ & ~new_n1380_ & ~new_n1397_ & new_n1381_;
  assign new_n1186_ = new_n1411_ & new_n1409_ & ~new_n1398_ & ~new_n1380_ & ~new_n1397_ & new_n1381_;
  assign new_n1187_ = new_n1411_ & ~new_n1409_ & ~new_n1398_ & ~new_n1380_ & ~new_n1397_ & new_n1381_;
  assign new_n1188_ = new_n1411_ & ~new_n1409_ & new_n1398_ & new_n1380_ & ~new_n1397_ & ~new_n1381_;
  assign new_n1189_ = new_n1411_ & ~new_n1409_ & ~new_n1398_ & new_n1380_ & ~new_n1397_ & ~new_n1381_;
  assign new_n1190_ = new_n1390_ & ~new_n1389_ & new_n1410_ & ~new_n1388_ & ~new_n1387_ & new_n1408_;
  assign new_n1191_ = ~new_n1411_ & ~new_n1409_ & new_n1398_ & new_n1380_ & ~new_n1397_ & ~new_n1381_;
  assign new_n1192_ = ~new_n1395_ & (pi198 ? pi019 : pi011);
  assign new_n1193_ = ~new_n1395_ & (pi198 ? pi020 : pi012);
  assign new_n1194_ = ~new_n1395_ & (pi198 ? pi021 : pi013);
  assign new_n1195_ = ~new_n1395_ & (pi198 ? pi022 : pi014);
  assign new_n1196_ = ~new_n1395_ & (pi198 ? pi023 : pi015);
  assign new_n1197_ = ~new_n1395_ & (pi198 ? pi024 : pi016);
  assign new_n1198_ = ~new_n1395_ & (pi198 ? pi025 : pi017);
  assign new_n1199_ = ~new_n1395_ & (pi198 ? pi026 : pi018);
  assign new_n1200_ = ~new_n1395_ & (pi198 ? pi027 : pi019);
  assign new_n1201_ = ~new_n1395_ & (pi198 ? pi028 : pi020);
  assign new_n1202_ = ~new_n1395_ & (pi198 ? pi029 : pi021);
  assign new_n1203_ = ~new_n1395_ & (pi198 ? pi030 : pi022);
  assign new_n1204_ = ~new_n1395_ & (pi198 ? pi031 : pi023);
  assign new_n1205_ = ~new_n1395_ & (pi198 ? pi032 : pi024);
  assign new_n1206_ = ~new_n1395_ & (pi198 ? pi033 : pi025);
  assign new_n1207_ = ~new_n1395_ & (pi198 ? pi034 : pi026);
  assign new_n1208_ = ~new_n1395_ & (pi198 ? pi035 : pi027);
  assign new_n1209_ = ~new_n1395_ & (pi198 ? pi036 : pi028);
  assign new_n1210_ = ~new_n1395_ & (pi198 ? pi037 : pi029);
  assign new_n1211_ = ~new_n1395_ & (pi198 ? pi038 : pi030);
  assign new_n1212_ = ~new_n1395_ & (pi198 ? pi039 : pi031);
  assign new_n1213_ = ~new_n1395_ & (pi198 ? pi040 : pi032);
  assign new_n1214_ = ~new_n1395_ & (pi198 ? pi041 : pi033);
  assign new_n1215_ = ~new_n1395_ & (pi198 ? pi042 : pi034);
  assign new_n1216_ = ~new_n1395_ & (pi198 ? pi043 : pi035);
  assign new_n1217_ = ~new_n1395_ & (pi198 ? pi044 : pi036);
  assign new_n1218_ = ~new_n1395_ & (pi198 ? pi045 : pi037);
  assign new_n1219_ = ~new_n1395_ & (pi198 ? pi046 : pi038);
  assign new_n1220_ = ~new_n1395_ & (pi198 ? pi047 : pi039);
  assign new_n1221_ = ~new_n1395_ & (pi198 ? pi048 : pi040);
  assign new_n1222_ = ~new_n1395_ & (pi198 ? pi049 : pi041);
  assign new_n1223_ = ~new_n1395_ & (pi198 ? pi050 : pi042);
  assign new_n1224_ = ~new_n1395_ & (pi198 ? pi051 : pi043);
  assign new_n1225_ = ~new_n1395_ & (pi198 ? pi052 : pi044);
  assign new_n1226_ = ~new_n1395_ & (pi198 ? pi053 : pi045);
  assign new_n1227_ = ~new_n1395_ & (pi198 ? pi054 : pi046);
  assign new_n1228_ = ~new_n1395_ & (pi198 ? pi055 : pi047);
  assign new_n1229_ = ~new_n1395_ & (pi198 ? pi056 : pi048);
  assign new_n1230_ = ~new_n1395_ & (pi198 ? pi057 : pi049);
  assign new_n1231_ = ~new_n1395_ & (pi198 ? pi058 : pi050);
  assign new_n1232_ = ~new_n1395_ & (pi198 ? pi059 : pi051);
  assign new_n1233_ = ~new_n1395_ & (pi198 ? pi060 : pi052);
  assign new_n1234_ = ~new_n1395_ & (pi198 ? pi061 : pi053);
  assign new_n1235_ = ~new_n1395_ & (pi198 ? pi062 : pi054);
  assign new_n1236_ = ~new_n1395_ & (pi198 ? pi063 : pi055);
  assign new_n1237_ = ~new_n1395_ & (pi198 ? pi064 : pi056);
  assign new_n1238_ = ~new_n1395_ & (pi198 ? pi065 : pi057);
  assign new_n1239_ = ~new_n1395_ & (pi198 ? pi066 : pi058);
  assign new_n1240_ = ~new_n1395_ & (pi198 ? pi000 : pi059);
  assign new_n1241_ = ~new_n1395_ & (pi198 ? pi001 : pi060);
  assign new_n1242_ = ~new_n1395_ & (pi198 ? pi002 : pi061);
  assign new_n1243_ = ~new_n1395_ & (pi198 ? pi003 : pi062);
  assign new_n1244_ = ~new_n1395_ & (pi198 ? pi004 : pi063);
  assign new_n1245_ = ~new_n1395_ & (pi198 ? pi005 : pi064);
  assign new_n1246_ = ~new_n1395_ & (pi198 ? pi006 : pi065);
  assign new_n1247_ = ~new_n1395_ & (pi198 ? pi007 : pi066);
  assign new_n1248_ = new_n1395_ ? pi017 : pi162;
  assign new_n1249_ = new_n1395_ ? pi025 : pi161;
  assign new_n1250_ = new_n1395_ ? pi033 : pi160;
  assign new_n1251_ = new_n1395_ ? pi041 : pi159;
  assign new_n1252_ = new_n1395_ ? pi049 : pi158;
  assign new_n1253_ = new_n1395_ ? pi057 : pi157;
  assign new_n1254_ = new_n1395_ ? pi065 : pi156;
  assign new_n1255_ = new_n1395_ ? pi006 : pi155;
  assign new_n1256_ = new_n1395_ ? pi015 : pi154;
  assign new_n1257_ = new_n1395_ ? pi023 : pi153;
  assign new_n1258_ = new_n1395_ ? pi031 : pi152;
  assign new_n1259_ = new_n1395_ ? pi039 : pi151;
  assign new_n1260_ = new_n1395_ ? pi047 : pi150;
  assign new_n1261_ = new_n1395_ ? pi055 : pi149;
  assign new_n1262_ = new_n1395_ ? pi063 : pi148;
  assign new_n1263_ = new_n1395_ ? pi004 : pi147;
  assign new_n1264_ = new_n1395_ ? pi013 : pi146;
  assign new_n1265_ = new_n1395_ ? pi021 : pi145;
  assign new_n1266_ = new_n1395_ ? pi029 : pi144;
  assign new_n1267_ = new_n1395_ ? pi037 : pi143;
  assign new_n1268_ = new_n1395_ ? pi045 : pi142;
  assign new_n1269_ = new_n1395_ ? pi053 : pi141;
  assign new_n1270_ = new_n1395_ ? pi061 : pi140;
  assign new_n1271_ = new_n1395_ ? pi002 : pi139;
  assign new_n1272_ = new_n1395_ ? pi011 : pi138;
  assign new_n1273_ = new_n1395_ ? pi019 : pi137;
  assign new_n1274_ = new_n1395_ ? pi027 : pi136;
  assign new_n1275_ = new_n1395_ ? pi035 : pi135;
  assign new_n1276_ = new_n1395_ ? pi043 : pi134;
  assign new_n1277_ = new_n1395_ ? pi051 : pi133;
  assign new_n1278_ = new_n1395_ ? pi059 : pi132;
  assign new_n1279_ = new_n1395_ ? pi000 : pi131;
  assign new_n1280_ = ~new_n1411_ & new_n1409_ & ~new_n1398_ & new_n1380_ & ~new_n1397_ & ~new_n1381_;
  assign new_n1281_ = ~new_n1411_ & ~new_n1409_ & new_n1398_ & ~new_n1380_ & ~new_n1397_ & ~new_n1381_;
  assign new_n1282_ = ~new_n1411_ & ~new_n1409_ & ~new_n1398_ & ~new_n1380_ & ~new_n1397_ & ~new_n1381_;
  assign new_n1283_ = ~new_n1394_ & new_n1393_ & ~new_n1414_ & ~new_n1392_ & ~new_n1412_ & new_n1391_;
  assign new_n1284_ = ~new_n1390_ & new_n1389_ & new_n1410_ & ~new_n1388_ & new_n1387_ & new_n1408_;
  assign new_n1285_ = new_n1395_ ? pi162 : (~pi198 & pi074);
  assign new_n1286_ = (pi255 & (~pi196 | ~pi195 | ~pi198 | ~pi197)) | (pi197 & pi196 & pi195 & pi009 & pi198);
  assign new_n1287_ = ~pi008 & (new_n1407_ ? (pi009 ? pi012 : pi004) : (new_n1403_ ? pi227 : (pi255 ? (new_n1405_ ? pi254 : pi253) : (new_n1405_ ? pi228 : pi229))));
  assign new_n1288_ = ~pi008 & (new_n1407_ ? (pi009 ? pi004 : pi063) : (new_n1403_ ? pi228 : (pi255 ? (new_n1405_ ? pi227 : pi254) : (new_n1405_ ? pi229 : pi230))));
  assign new_n1289_ = ~pi008 & (new_n1407_ ? (pi009 ? pi063 : pi055) : (new_n1403_ ? pi229 : (pi255 ? (new_n1405_ ? pi228 : pi227) : (new_n1405_ ? pi230 : pi231))));
  assign new_n1290_ = ~pi008 & (new_n1407_ ? (pi009 ? pi055 : pi047) : (new_n1403_ ? pi230 : (pi255 ? (new_n1405_ ? pi229 : pi228) : (new_n1405_ ? pi231 : pi232))));
  assign new_n1291_ = ~pi008 & (new_n1407_ ? (pi009 ? pi047 : pi003) : (new_n1403_ ? pi231 : (pi255 ? (new_n1405_ ? pi230 : pi229) : (new_n1405_ ? pi232 : pi233))));
  assign new_n1292_ = ~pi008 & (new_n1407_ ? (pi009 ? pi003 : pi062) : (new_n1403_ ? pi232 : (pi255 ? (new_n1405_ ? pi231 : pi230) : (new_n1405_ ? pi233 : pi234))));
  assign new_n1293_ = ~pi008 & (new_n1407_ ? (pi009 ? pi062 : pi054) : (new_n1403_ ? pi233 : (pi255 ? (new_n1405_ ? pi232 : pi231) : (new_n1405_ ? pi234 : pi235))));
  assign new_n1294_ = new_n1395_ ? pi145 : (pi198 ? pi070 : pi078);
  assign new_n1295_ = ~pi008 & (new_n1407_ ? (pi009 ? pi046 : pi038) : (new_n1403_ ? pi235 : (pi255 ? (new_n1405_ ? pi234 : pi233) : (new_n1405_ ? pi236 : pi237))));
  assign new_n1296_ = ~pi008 & (new_n1407_ ? (pi009 ? pi038 : pi030) : (new_n1403_ ? pi236 : (pi255 ? (new_n1405_ ? pi235 : pi234) : (new_n1405_ ? pi237 : pi238))));
  assign new_n1297_ = ~pi008 & (new_n1407_ ? (pi009 ? pi030 : pi022) : (new_n1403_ ? pi237 : (pi255 ? (new_n1405_ ? pi236 : pi235) : (new_n1405_ ? pi238 : pi239))));
  assign new_n1298_ = ~pi008 & (new_n1407_ ? (pi009 ? pi022 : pi014) : (new_n1403_ ? pi238 : (pi255 ? (new_n1405_ ? pi237 : pi236) : (new_n1405_ ? pi239 : pi240))));
  assign new_n1299_ = ~pi008 & (new_n1407_ ? (pi009 ? pi014 : pi002) : (new_n1403_ ? pi239 : (pi255 ? (new_n1405_ ? pi238 : pi237) : (new_n1405_ ? pi240 : pi241))));
  assign new_n1300_ = ~pi008 & (new_n1407_ ? (pi009 ? pi002 : pi061) : (new_n1403_ ? pi240 : (pi255 ? (new_n1405_ ? pi239 : pi238) : (new_n1405_ ? pi241 : pi242))));
  assign new_n1301_ = ~pi008 & (new_n1407_ ? (pi009 ? pi061 : pi053) : (new_n1403_ ? pi241 : (pi255 ? (new_n1405_ ? pi240 : pi239) : (new_n1405_ ? pi242 : pi243))));
  assign new_n1302_ = ~pi008 & (new_n1407_ ? (pi009 ? pi053 : pi045) : (new_n1403_ ? pi242 : (pi255 ? (new_n1405_ ? pi241 : pi240) : (new_n1405_ ? pi243 : pi244))));
  assign new_n1303_ = ~pi008 & (new_n1407_ ? (pi009 ? pi045 : pi037) : (new_n1403_ ? pi243 : (pi255 ? (new_n1405_ ? pi242 : pi241) : (new_n1405_ ? pi244 : pi245))));
  assign new_n1304_ = ~pi008 & (new_n1407_ ? (pi009 ? pi037 : pi029) : (new_n1403_ ? pi244 : (pi255 ? (new_n1405_ ? pi243 : pi242) : (new_n1405_ ? pi245 : pi246))));
  assign new_n1305_ = ~pi008 & (new_n1407_ ? (pi009 ? pi029 : pi021) : (new_n1403_ ? pi245 : (pi255 ? (new_n1405_ ? pi244 : pi243) : (new_n1405_ ? pi246 : pi247))));
  assign new_n1306_ = ~pi008 & (new_n1407_ ? (pi009 ? pi021 : pi013) : (new_n1403_ ? pi246 : (pi255 ? (new_n1405_ ? pi245 : pi244) : (new_n1405_ ? pi247 : pi248))));
  assign new_n1307_ = new_n1395_ ? pi155 : (pi198 ? pi122 : pi130);
  assign new_n1308_ = ~pi008 & (new_n1407_ ? (pi009 ? pi054 : pi046) : (new_n1403_ ? pi234 : (pi255 ? (new_n1405_ ? pi233 : pi232) : (new_n1405_ ? pi235 : pi236))));
  assign new_n1309_ = new_n1395_ ? pi147 : (pi198 ? pi120 : pi128);
  assign new_n1310_ = new_n1395_ ? pi154 : (~pi198 & pi072);
  assign new_n1311_ = new_n1395_ ? pi139 : (pi198 ? pi118 : pi126);
  assign new_n1312_ = ~pi008 & (new_n1407_ ? (pi009 ? pi001 : pi060) : (new_n1403_ ? pi248 : (pi255 ? (new_n1405_ ? pi247 : pi246) : (new_n1405_ ? pi249 : pi250))));
  assign new_n1313_ = new_n1395_ ? pi131 : (pi198 ? pi116 : pi124);
  assign new_n1314_ = ~pi008 & (new_n1407_ ? (pi009 ? pi013 : pi001) : (new_n1403_ ? pi247 : (pi255 ? (new_n1405_ ? pi246 : pi245) : (new_n1405_ ? pi248 : pi249))));
  assign new_n1315_ = new_n1395_ ? pi156 : (pi198 ? pi114 : pi122);
  assign new_n1316_ = new_n1395_ ? pi146 : (~pi198 & pi070);
  assign new_n1317_ = new_n1395_ ? pi148 : (pi198 ? pi112 : pi120);
  assign new_n1318_ = ~pi008 & (new_n1407_ ? (pi009 ? pi052 : pi044) : (new_n1403_ ? pi250 : (pi255 ? (new_n1405_ ? pi249 : pi248) : (new_n1405_ ? pi251 : pi252))));
  assign new_n1319_ = new_n1395_ ? pi140 : (pi198 ? pi110 : pi118);
  assign new_n1320_ = ~pi008 & (new_n1407_ ? (pi009 ? pi060 : pi052) : (new_n1403_ ? pi249 : (pi255 ? (new_n1405_ ? pi248 : pi247) : (new_n1405_ ? pi250 : pi251))));
  assign new_n1321_ = new_n1395_ ? pi132 : (pi198 ? pi108 : pi116);
  assign new_n1322_ = new_n1395_ ? pi138 : (~pi198 & pi068);
  assign new_n1323_ = new_n1395_ ? pi157 : (pi198 ? pi106 : pi114);
  assign new_n1324_ = ~pi008 & (new_n1407_ ? (pi009 ? pi036 : pi028) : (new_n1403_ ? pi252 : (pi255 ? (new_n1405_ ? pi251 : pi250) : (new_n1405_ ? pi253 : pi254))));
  assign new_n1325_ = new_n1395_ ? pi149 : (pi198 ? pi104 : pi112);
  assign new_n1326_ = ~pi008 & (new_n1407_ ? (pi009 ? pi044 : pi036) : (new_n1403_ ? pi251 : (pi255 ? (new_n1405_ ? pi250 : pi249) : (new_n1405_ ? pi252 : pi253))));
  assign new_n1327_ = new_n1395_ ? pi141 : (pi198 ? pi102 : pi110);
  assign new_n1328_ = ~pi008 & (new_n1407_ ? (pi009 ? pi020 : pi012) : (new_n1403_ ? pi254 : (pi255 ? (new_n1405_ ? pi253 : pi252) : (new_n1405_ ? pi227 : pi228))));
  assign new_n1329_ = new_n1395_ ? pi133 : (pi198 ? pi100 : pi108);
  assign new_n1330_ = ~pi008 & (new_n1407_ ? (pi009 ? pi028 : pi020) : (new_n1403_ ? pi253 : (pi255 ? (new_n1405_ ? pi252 : pi251) : (new_n1405_ ? pi254 : pi227))));
  assign new_n1331_ = new_n1395_ ? pi158 : (pi198 ? pi098 : pi106);
  assign new_n1332_ = ~pi008 & (new_n1407_ ? (pi009 ? pi039 : pi031) : (new_n1403_ ? pi200 : (pi255 ? (new_n1405_ ? pi199 : pi226) : (new_n1405_ ? pi201 : pi202))));
  assign new_n1333_ = new_n1395_ ? pi150 : (pi198 ? pi096 : pi104);
  assign new_n1334_ = ~pi008 & (new_n1407_ ? (pi009 ? pi018 : pi039) : (new_n1403_ ? pi199 : (pi255 ? (new_n1405_ ? pi226 : pi225) : (new_n1405_ ? pi200 : pi201))));
  assign new_n1335_ = new_n1395_ ? pi142 : (pi198 ? pi094 : pi102);
  assign new_n1336_ = ~pi008 & (new_n1407_ ? (pi009 ? pi023 : pi015) : (new_n1403_ ? pi202 : (pi255 ? (new_n1405_ ? pi201 : pi200) : (new_n1405_ ? pi203 : pi204))));
  assign new_n1337_ = new_n1395_ ? pi134 : (pi198 ? pi092 : pi100);
  assign new_n1338_ = ~pi008 & (new_n1407_ ? (pi009 ? pi031 : pi023) : (new_n1403_ ? pi201 : (pi255 ? (new_n1405_ ? pi200 : pi199) : (new_n1405_ ? pi202 : pi203))));
  assign new_n1339_ = new_n1395_ ? pi159 : (pi198 ? pi090 : pi098);
  assign new_n1340_ = ~pi008 & (new_n1407_ ? (pi009 ? pi005 : pi064) : (new_n1403_ ? pi204 : (pi255 ? (new_n1405_ ? pi203 : pi202) : (new_n1405_ ? pi205 : pi206))));
  assign new_n1341_ = new_n1395_ ? pi151 : (pi198 ? pi088 : pi096);
  assign new_n1342_ = ~pi008 & (new_n1407_ ? (pi009 ? pi015 : pi005) : (new_n1403_ ? pi203 : (pi255 ? (new_n1405_ ? pi202 : pi201) : (new_n1405_ ? pi204 : pi205))));
  assign new_n1343_ = new_n1395_ ? pi143 : (pi198 ? pi086 : pi094);
  assign new_n1344_ = ~pi008 & (new_n1407_ ? (pi009 ? pi056 : pi048) : (new_n1403_ ? pi206 : (pi255 ? (new_n1405_ ? pi205 : pi204) : (new_n1405_ ? pi207 : pi208))));
  assign new_n1345_ = new_n1395_ ? pi135 : (pi198 ? pi084 : pi092);
  assign new_n1346_ = ~pi008 & (new_n1407_ ? (pi009 ? pi064 : pi056) : (new_n1403_ ? pi205 : (pi255 ? (new_n1405_ ? pi204 : pi203) : (new_n1405_ ? pi206 : pi207))));
  assign new_n1347_ = new_n1395_ ? pi160 : (pi198 ? pi082 : pi090);
  assign new_n1348_ = ~pi008 & (new_n1407_ ? (pi009 ? pi040 : pi032) : (new_n1403_ ? pi208 : (pi255 ? (new_n1405_ ? pi207 : pi206) : (new_n1405_ ? pi209 : pi210))));
  assign new_n1349_ = new_n1395_ ? pi152 : (pi198 ? pi080 : pi088);
  assign new_n1350_ = ~pi008 & (new_n1407_ ? (pi009 ? pi048 : pi040) : (new_n1403_ ? pi207 : (pi255 ? (new_n1405_ ? pi206 : pi205) : (new_n1405_ ? pi208 : pi209))));
  assign new_n1351_ = new_n1395_ ? pi144 : (pi198 ? pi078 : pi086);
  assign new_n1352_ = new_n1395_ ? pi136 : (pi198 ? pi076 : pi084);
  assign new_n1353_ = new_n1395_ ? pi161 : (pi198 ? pi074 : pi082);
  assign new_n1354_ = ~pi008 & (new_n1407_ ? (pi009 ? pi024 : pi016) : (new_n1403_ ? pi210 : (pi255 ? (new_n1405_ ? pi209 : pi208) : (new_n1405_ ? pi211 : pi212))));
  assign new_n1355_ = new_n1395_ ? pi153 : (pi198 ? pi072 : pi080);
  assign new_n1356_ = ~pi008 & (new_n1407_ ? (pi009 ? pi032 : pi024) : (new_n1403_ ? pi209 : (pi255 ? (new_n1405_ ? pi208 : pi207) : (new_n1405_ ? pi210 : pi211))));
  assign new_n1357_ = ~pi008 & (new_n1407_ ? (pi009 ? pi016 : pi006) : (new_n1403_ ? pi211 : (pi255 ? (new_n1405_ ? pi210 : pi209) : (new_n1405_ ? pi212 : pi213))));
  assign new_n1358_ = ~pi008 & (new_n1407_ ? (pi009 ? pi006 : pi065) : (new_n1403_ ? pi212 : (pi255 ? (new_n1405_ ? pi211 : pi210) : (new_n1405_ ? pi213 : pi214))));
  assign new_n1359_ = new_n1395_ ? pi137 : (pi198 ? pi068 : pi076);
  assign new_n1360_ = ~pi198 & ~new_n1407_ & ~pi008;
  assign new_n1361_ = ~pi008 & (new_n1407_ ? (pi009 ? pi065 : pi057) : (new_n1403_ ? pi213 : (pi255 ? (new_n1405_ ? pi212 : pi211) : (new_n1405_ ? pi214 : pi215))));
  assign new_n1362_ = ~pi008 & (new_n1407_ ? (pi009 ? pi057 : pi049) : (new_n1403_ ? pi214 : (pi255 ? (new_n1405_ ? pi213 : pi212) : (new_n1405_ ? pi215 : pi216))));
  assign new_n1363_ = ~pi008 & (new_n1407_ ? (pi009 ? pi049 : pi041) : (new_n1403_ ? pi215 : (pi255 ? (new_n1405_ ? pi214 : pi213) : (new_n1405_ ? pi216 : pi217))));
  assign new_n1364_ = ~pi008 & (new_n1407_ ? (pi009 ? pi041 : pi033) : (new_n1403_ ? pi216 : (pi255 ? (new_n1405_ ? pi215 : pi214) : (new_n1405_ ? pi217 : pi218))));
  assign new_n1365_ = ~pi008 & (new_n1407_ ? (pi009 ? pi033 : pi025) : (new_n1403_ ? pi217 : (pi255 ? (new_n1405_ ? pi216 : pi215) : (new_n1405_ ? pi218 : pi219))));
  assign new_n1366_ = ~pi008 & (new_n1407_ ? (pi009 ? pi025 : pi017) : (new_n1403_ ? pi218 : (pi255 ? (new_n1405_ ? pi217 : pi216) : (new_n1405_ ? pi219 : pi220))));
  assign new_n1367_ = ~pi008 & (new_n1407_ ? (pi009 ? pi017 : pi007) : (new_n1403_ ? pi219 : (pi255 ? (new_n1405_ ? pi218 : pi217) : (new_n1405_ ? pi220 : pi221))));
  assign new_n1368_ = ~pi008 & (new_n1407_ ? (pi009 ? pi007 : pi066) : (new_n1403_ ? pi220 : (pi255 ? (new_n1405_ ? pi219 : pi218) : (new_n1405_ ? pi221 : pi222))));
  assign new_n1369_ = ~pi008 & (new_n1407_ ? (pi009 ? pi066 : pi058) : (new_n1403_ ? pi221 : (pi255 ? (new_n1405_ ? pi220 : pi219) : (new_n1405_ ? pi222 : pi223))));
  assign new_n1370_ = ~pi008 & (new_n1407_ ? (pi009 ? pi058 : pi050) : (new_n1403_ ? pi222 : (pi255 ? (new_n1405_ ? pi221 : pi220) : (new_n1405_ ? pi223 : pi224))));
  assign new_n1371_ = ~pi008 & (new_n1407_ ? (pi009 ? pi050 : pi042) : (new_n1403_ ? pi223 : (pi255 ? (new_n1405_ ? pi222 : pi221) : (new_n1405_ ? pi224 : pi225))));
  assign new_n1372_ = ~pi008 & (new_n1407_ ? (pi009 ? pi042 : pi034) : (new_n1403_ ? pi224 : (pi255 ? (new_n1405_ ? pi223 : pi222) : (new_n1405_ ? pi225 : pi226))));
  assign new_n1373_ = ~pi008 & (new_n1407_ ? (pi009 ? pi034 : pi026) : (new_n1403_ ? pi225 : (pi255 ? (new_n1405_ ? pi224 : pi223) : (new_n1405_ ? pi226 : pi199))));
  assign new_n1374_ = ~pi008 & (new_n1407_ ? (pi009 ? pi026 : pi018) : (new_n1403_ ? pi226 : (pi255 ? (new_n1405_ ? pi225 : pi224) : (new_n1405_ ? pi199 : pi200))));
  assign new_n1375_ = ~new_n1407_ & ~pi008 & (pi198 ^ pi197);
  assign new_n1376_ = pi208 ^ pi154;
  assign new_n1377_ = pi206 ^ pi155;
  assign new_n1378_ = pi204 ^ pi155;
  assign new_n1379_ = pi212 ^ pi157;
  assign new_n1380_ = pi216 ^ pi161;
  assign new_n1381_ = pi210 ^ pi162;
  assign new_n1382_ = pi215 ^ pi153;
  assign new_n1383_ = pi201 ^ pi151;
  assign new_n1384_ = pi211 ^ pi151;
  assign new_n1385_ = pi200 ^ pi149;
  assign new_n1386_ = pi214 ^ pi147;
  assign new_n1387_ = pi242 ^ pi147;
  assign new_n1388_ = pi252 ^ pi145;
  assign new_n1389_ = pi236 ^ pi143;
  assign new_n1390_ = pi228 ^ pi142;
  assign new_n1391_ = pi243 ^ pi142;
  assign new_n1392_ = pi232 ^ pi141;
  assign new_n1393_ = pi250 ^ pi139;
  assign new_n1394_ = pi235 ^ pi138;
  assign new_n1395_ = pi195 & pi196 & pi198 & pi197;
  assign new_n1396_ = pi221 ^ pi156;
  assign new_n1397_ = pi213 ^ pi131;
  assign new_n1398_ = pi203 ^ pi160;
  assign new_n1399_ = pi217 ^ pi154;
  assign new_n1400_ = pi223 ^ pi152;
  assign new_n1401_ = pi219 ^ pi150;
  assign new_n1402_ = pi220 ^ pi150;
  assign new_n1403_ = pi198 & pi197 & pi196 & pi195 & (pi009 ^ pi255);
  assign new_n1404_ = pi207 ^ pi148;
  assign new_n1405_ = (pi197 & pi196 & (pi198 | (~pi198 & pi195))) | (~pi198 & ~pi197 & ~pi196 & ~pi195);
  assign new_n1406_ = pi225 ^ pi146;
  assign new_n1407_ = pi010 & pi195 & pi196 & pi198 & pi197;
  assign new_n1408_ = pi231 ^ pi146;
  assign new_n1409_ = pi226 ^ pi159;
  assign new_n1410_ = pi246 ^ pi144;
  assign new_n1411_ = pi222 ^ pi158;
  assign new_n1412_ = pi253 ^ pi143;
  assign new_n1413_ = pi224 ^ pi159;
  assign new_n1414_ = pi238 ^ pi140;
  assign new_n1415_ = pi239 ^ pi139;
  assign new_n1416_ = pi234 ^ pi138;
  assign new_n1417_ = pi244 ^ pi137;
  assign new_n1418_ = pi227 ^ pi136;
  assign new_n1419_ = pi249 ^ pi135;
  assign new_n1420_ = pi230 ^ pi134;
  assign new_n1421_ = pi237 ^ pi135;
  assign new_n1422_ = pi241 ^ pi134;
  assign new_n1423_ = pi233 ^ pi133;
  assign new_n1424_ = pi247 ^ pi132;
  assign new_n1425_ = pi254 ^ pi131;
  assign new_n1426_ = pi251 ^ pi162;
  assign new_n1427_ = pi199 ^ pi158;
endmodule


