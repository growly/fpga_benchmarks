// Benchmark "k2" written by ABC on Thu Mar 19 13:02:36 2020

module k2 ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44;
  wire new_n116_, new_n135_, new_n136_, new_n137_, new_n138_, new_n139_,
    new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_,
    new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_,
    new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_,
    new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_,
    new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_,
    new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_,
    new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_,
    new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_,
    new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_,
    new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_,
    new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_,
    new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_,
    new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_,
    new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_,
    new_n314_, new_n315_;
  assign po00 = new_n279_ | new_n229_ | new_n246_ | new_n228_ | new_n222_ | new_n149_;
  assign po01 = new_n222_ | new_n279_;
  assign po03 = new_n228_ | new_n229_;
  assign po04 = new_n279_ | new_n149_ | new_n229_;
  assign po05 = new_n223_ | new_n150_ | new_n247_ | new_n261_;
  assign po06 = new_n196_ | new_n203_ | new_n199_ | new_n138_ | new_n137_ | new_n142_ | new_n139_ | new_n148_ | new_n153_ | new_n154_ | new_n156_ | new_n158_ | new_n310_ | new_n315_ | new_n286_ | new_n304_ | new_n291_ | new_n297_ | new_n273_ | new_n287_ | new_n267_ | new_n270_ | new_n212_ | new_n216_ | new_n217_ | new_n218_ | new_n252_ | new_n264_ | new_n219_ | po41;
  assign po07 = new_n142_ | new_n267_ | new_n153_ | new_n264_ | new_n216_ | new_n217_;
  assign po08 = new_n199_ | new_n142_ | new_n137_ | new_n156_ | new_n148_ | new_n304_ | new_n286_ | new_n212_ | new_n216_ | new_n218_ | po41 | new_n270_ | new_n287_ | new_n252_ | new_n264_;
  assign po09 = new_n196_ | new_n291_ | new_n297_;
  assign po10 = new_n183_ | new_n180_ | new_n184_ | new_n186_ | new_n185_ | new_n187_ | new_n189_ | new_n188_ | new_n193_ | new_n198_ | new_n195_ | new_n136_ | new_n202_ | new_n143_ | new_n147_ | new_n144_ | po21 | new_n300_ | po20 | new_n285_ | new_n302_ | new_n314_ | new_n305_ | new_n307_ | new_n167_ | new_n288_ | new_n292_ | new_n239_ | new_n274_ | new_n275_ | new_n272_ | new_n268_ | new_n271_ | new_n231_ | new_n224_ | new_n230_ | new_n221_ | new_n213_ | new_n220_ | new_n253_ | new_n265_ | new_n248_ | new_n152_ | new_n240_;
  assign po11 = new_n195_ | new_n178_ | new_n202_ | new_n197_ | new_n143_ | new_n141_ | new_n155_ | new_n314_ | new_n300_ | new_n167_ | new_n305_ | new_n292_ | new_n239_ | new_n288_ | new_n274_ | new_n275_ | new_n272_ | new_n269_ | new_n271_ | new_n265_ | new_n266_ | new_n254_ | new_n249_ | new_n253_ | new_n241_ | new_n248_ | new_n240_ | new_n152_ | new_n157_ | new_n233_ | new_n234_ | new_n231_ | new_n225_ | new_n230_ | new_n221_ | new_n224_ | new_n220_ | new_n213_ | new_n214_;
  assign po12 = new_n179_ | new_n193_ | new_n180_ | new_n195_ | new_n198_ | new_n197_ | new_n202_ | new_n141_ | new_n136_ | po21 | new_n147_ | new_n144_ | new_n143_ | po20 | new_n300_ | new_n155_ | new_n285_ | new_n302_ | new_n314_ | new_n307_ | new_n167_ | new_n305_ | new_n288_ | new_n292_ | new_n239_ | new_n243_ | new_n274_ | new_n271_ | new_n272_ | new_n235_ | new_n275_ | new_n227_ | new_n269_ | new_n266_ | new_n268_ | new_n254_ | new_n265_ | new_n249_ | new_n253_ | new_n248_ | new_n240_ | new_n241_ | new_n157_ | new_n234_ | new_n152_ | new_n213_ | new_n214_ | new_n220_ | new_n221_ | new_n233_ | new_n224_ | new_n225_;
  assign po13 = new_n162_ | new_n161_ | new_n282_ | new_n308_ | new_n285_ | new_n312_ | new_n303_ | new_n309_ | new_n302_ | new_n307_ | new_n263_ | new_n227_ | new_n231_ | new_n268_ | new_n230_ | new_n207_ | new_n210_ | new_n296_ | new_n306_ | new_n283_ | new_n235_ | new_n243_ | new_n140_ | new_n141_ | new_n144_ | new_n147_ | new_n145_ | new_n151_ | po20 | po21 | new_n155_ | new_n160_ | new_n159_ | new_n183_ | new_n180_ | new_n184_ | new_n186_ | new_n185_ | new_n197_ | new_n189_ | new_n198_ | new_n136_ | new_n298_;
  assign po14 = new_n181_ | new_n185_ | new_n183_ | new_n189_ | new_n187_ | new_n197_ | new_n192_ | new_n198_ | new_n141_ | new_n136_ | po20 | po21 | new_n147_ | new_n144_ | new_n221_ | new_n231_ | new_n157_ | new_n241_ | new_n275_ | new_n268_ | new_n272_ | new_n155_ | new_n285_ | new_n282_ | new_n302_ | new_n308_ | new_n235_ | new_n307_;
  assign po15 = new_n306_ | new_n304_ | new_n305_ | new_n284_ | new_n299_ | new_n293_ | new_n167_ | new_n291_ | new_n292_ | new_n245_ | new_n288_ | new_n239_ | new_n244_ | new_n271_ | new_n274_ | new_n268_ | new_n253_ | new_n265_ | new_n248_ | new_n250_ | new_n240_ | new_n247_ | new_n207_ | new_n210_ | new_n213_ | new_n220_ | new_n231_ | new_n152_ | new_n224_ | new_n230_ | new_n170_ | new_n173_ | new_n172_ | new_n176_ | new_n175_ | new_n178_ | new_n177_ | new_n196_ | new_n195_ | new_n194_ | new_n182_ | new_n200_ | new_n198_ | new_n204_ | new_n202_ | new_n136_ | new_n140_ | new_n143_ | po20 | po21 | new_n147_ | new_n144_ | new_n160_ | new_n300_ | new_n285_ | new_n236_ | new_n307_ | new_n302_ | new_n313_ | new_n314_;
  assign po16 = new_n180_ | new_n184_ | new_n183_ | new_n185_ | new_n187_ | new_n186_ | new_n188_ | new_n193_ | new_n189_ | new_n196_ | new_n194_ | new_n198_ | new_n197_ | new_n200_ | new_n204_ | new_n202_ | new_n298_ | new_n206_ | new_n141_ | new_n136_ | new_n140_ | new_n145_ | new_n144_ | po20 | po21 | new_n151_ | new_n147_ | new_n207_ | new_n210_ | new_n220_ | new_n268_ | new_n244_ | new_n271_ | new_n274_ | new_n304_ | new_n284_ | new_n299_ | new_n116_ | new_n294_ | new_n245_ | new_n291_ | new_n285_ | new_n313_ | new_n308_ | new_n307_ | new_n302_ | new_n309_ | new_n312_ | new_n155_ | new_n160_ | new_n159_ | new_n162_ | new_n282_ | new_n236_;
  assign po17 = new_n171_ | new_n170_ | new_n178_ | new_n177_ | new_n181_ | new_n179_ | new_n192_ | new_n182_ | new_n195_ | new_n194_ | new_n206_ | new_n198_ | new_n143_ | new_n144_ | new_n140_ | new_n141_ | new_n136_ | po21 | new_n147_ | new_n155_ | po20 | new_n162_ | new_n161_ | new_n160_ | new_n300_ | new_n314_ | new_n308_ | new_n285_ | new_n282_ | new_n306_ | new_n309_ | new_n305_ | new_n293_ | new_n167_ | new_n227_ | new_n235_ | new_n275_ | new_n276_ | new_n239_ | new_n243_ | new_n288_ | new_n292_ | new_n254_ | new_n265_ | new_n253_ | new_n249_ | new_n251_ | new_n266_ | new_n268_ | new_n269_ | new_n272_ | new_n241_ | new_n248_ | new_n157_ | new_n240_ | new_n234_ | new_n152_ | new_n231_ | new_n233_ | new_n214_ | new_n220_ | new_n213_ | new_n207_ | new_n210_ | new_n221_ | new_n224_ | new_n225_ | new_n230_;
  assign po18 = new_n171_ | new_n170_ | new_n172_ | new_n194_ | new_n173_ | new_n195_ | new_n298_ | new_n197_ | new_n143_ | new_n151_ | new_n145_ | new_n159_ | new_n300_ | new_n162_ | new_n314_ | new_n165_ | new_n312_ | new_n303_ | new_n309_ | new_n302_ | new_n307_ | new_n263_ | new_n305_ | new_n306_ | new_n167_ | new_n293_ | new_n296_ | new_n292_ | new_n283_ | new_n288_ | new_n239_ | new_n253_ | new_n265_ | new_n231_ | new_n224_ | new_n230_ | new_n213_ | new_n207_ | new_n210_ | new_n248_ | new_n251_ | new_n247_ | new_n152_ | new_n240_;
  assign po19 = new_n172_ | new_n175_ | new_n174_ | new_n178_ | new_n194_ | new_n182_ | new_n298_ | new_n143_ | new_n141_ | new_n195_ | new_n202_ | new_n197_ | new_n140_ | new_n151_ | new_n145_ | new_n155_ | new_n159_ | new_n300_ | new_n160_ | new_n282_ | new_n161_ | new_n314_ | new_n308_ | new_n303_ | new_n309_ | new_n274_ | new_n265_ | new_n271_ | new_n253_ | new_n247_ | new_n248_ | new_n213_ | new_n220_ | new_n224_ | new_n230_ | new_n240_ | new_n231_ | new_n152_ | new_n302_ | new_n306_ | new_n263_ | new_n305_ | new_n296_ | new_n167_ | new_n294_ | new_n292_ | new_n116_ | new_n288_ | new_n239_ | new_n283_;
  assign po20 = pi30 & pi29 & ~pi28 & pi26 & ~pi21 & pi20 & ~pi19 & ~pi17 & pi18;
  assign po21 = ~pi30 & pi29 & pi28 & pi26 & ~pi21 & pi20 & pi18 & ~pi19;
  assign po22 = new_n170_ | new_n172_ | new_n171_ | new_n174_ | new_n173_ | new_n176_ | new_n175_ | new_n177_ | new_n179_ | new_n178_ | new_n181_ | new_n180_ | new_n183_ | new_n182_ | new_n184_ | new_n186_ | new_n185_ | new_n188_ | new_n187_ | new_n192_ | new_n189_ | new_n194_ | new_n193_ | new_n196_ | new_n195_ | new_n198_ | new_n197_ | new_n202_ | new_n200_ | new_n204_ | new_n298_ | new_n206_ | new_n141_ | new_n136_ | new_n140_ | new_n143_ | new_n144_ | new_n146_ | new_n145_ | new_n151_ | new_n147_ | po20 | po21 | new_n155_ | new_n159_ | new_n300_ | new_n161_ | new_n160_ | new_n163_ | new_n162_ | new_n236_ | new_n165_ | new_n285_ | new_n282_ | new_n314_ | new_n308_ | new_n312_ | new_n313_ | new_n269_ | new_n266_ | new_n268_ | new_n260_ | new_n265_ | new_n254_ | new_n259_ | new_n251_ | new_n253_ | new_n249_ | new_n250_ | new_n247_ | new_n248_ | new_n240_ | new_n241_ | new_n157_ | new_n234_ | new_n152_ | new_n232_ | new_n233_ | new_n230_ | new_n231_ | new_n207_ | new_n213_ | new_n214_ | new_n215_ | new_n224_ | new_n225_ | new_n220_ | new_n221_ | new_n291_ | new_n245_ | new_n288_ | new_n239_ | new_n243_ | new_n283_ | new_n244_ | new_n235_ | new_n278_ | new_n276_ | new_n227_ | new_n271_ | new_n272_ | new_n274_ | new_n275_ | new_n309_ | new_n302_ | new_n303_ | new_n307_ | new_n263_ | new_n304_ | new_n306_ | new_n299_ | new_n167_ | new_n284_ | new_n294_ | new_n296_ | new_n116_ | new_n293_;
  assign po23 = new_n274_ | new_n220_ | new_n271_;
  assign new_n116_ = pi30 & ~pi29 & pi22 & ~pi21 & pi20 & ~pi18 & ~pi19;
  assign po25 = new_n177_ | new_n140_ | new_n298_ | new_n146_ | new_n145_ | new_n159_ | new_n151_ | new_n161_ | new_n160_ | new_n163_ | new_n162_ | new_n258_ | new_n165_ | new_n309_ | new_n312_ | new_n303_ | new_n306_ | new_n263_ | new_n295_ | new_n296_ | new_n116_ | new_n293_ | new_n210_ | new_n215_ | new_n232_ | new_n259_ | new_n280_ | new_n283_ | new_n260_ | new_n278_;
  assign po26 = new_n283_ | new_n296_ | new_n303_ | new_n298_;
  assign po27 = new_n304_ | new_n284_ | new_n299_ | new_n291_ | new_n244_ | new_n245_ | new_n200_ | new_n196_ | new_n204_ | new_n313_ | new_n236_;
  assign po28 = new_n170_ | new_n169_ | new_n171_ | new_n173_ | new_n172_ | new_n175_ | new_n174_ | new_n176_ | new_n182_ | new_n179_ | new_n116_ | new_n280_ | new_n243_ | new_n278_ | new_n227_ | new_n235_ | new_n258_ | new_n294_ | new_n295_ | new_n165_ | new_n163_ | new_n233_ | new_n225_ | new_n232_ | new_n221_ | new_n214_ | new_n215_ | new_n164_ | new_n226_ | new_n237_ | new_n234_ | new_n157_ | new_n275_ | new_n276_ | new_n269_ | new_n168_ | new_n262_ | new_n259_ | new_n260_ | new_n135_ | new_n251_ | new_n257_;
  assign po29 = new_n158_ | new_n304_ | new_n315_ | new_n196_ | new_n139_ | new_n203_ | new_n261_ | new_n270_ | new_n273_ | new_n297_ | new_n287_ | new_n291_ | new_n223_ | new_n218_ | new_n219_ | new_n217_ | new_n212_ | new_n216_ | new_n247_ | new_n150_ | po41 | new_n267_ | new_n252_ | new_n264_;
  assign po30 = new_n199_ | new_n153_ | new_n142_ | new_n148_ | new_n286_ | new_n310_;
  assign po31 = new_n199_ | new_n138_ | new_n137_ | new_n156_ | new_n286_ | new_n154_;
  assign po32 = ~pi30 & ~pi29 & ~pi28 & ~pi27 & pi21 & ~pi14 & ~pi12 & ~pi13;
  assign po33 = new_n196_ | new_n195_ | new_n198_ | new_n204_ | new_n200_;
  assign po34 = new_n180_ | new_n178_ | new_n181_ | new_n185_ | new_n183_ | new_n186_ | new_n188_ | new_n187_ | new_n189_ | new_n191_ | new_n190_ | new_n192_ | new_n201_ | new_n199_ | new_n202_ | new_n137_ | new_n203_ | new_n156_ | new_n155_ | new_n154_ | new_n138_ | new_n143_ | new_n141_ | new_n241_ | new_n150_ | new_n152_ | new_n229_ | new_n149_ | new_n228_ | new_n254_ | new_n249_ | new_n250_ | new_n288_ | new_n266_ | new_n272_ | new_n167_ | new_n289_ | new_n291_ | new_n314_ | new_n277_ | new_n304_ | new_n282_ | new_n300_ | new_n286_ | new_n311_ | new_n308_;
  assign po35 = new_n184_ | new_n177_ | new_n195_ | new_n193_ | new_n199_ | new_n197_ | new_n200_ | new_n204_ | new_n201_ | new_n298_ | new_n206_ | new_n138_ | new_n137_ | new_n140_ | new_n139_ | new_n142_ | new_n145_ | new_n153_ | new_n151_ | new_n148_ | new_n154_ | new_n156_ | new_n158_ | new_n310_ | new_n159_ | new_n282_ | new_n160_ | new_n263_ | new_n303_ | new_n306_ | new_n281_ | new_n304_ | new_n315_ | new_n308_ | new_n286_ | new_n285_ | new_n290_ | new_n291_ | new_n287_ | new_n239_ | new_n283_ | new_n293_ | new_n296_ | new_n297_ | new_n301_ | new_n274_ | new_n261_ | new_n271_ | new_n273_ | new_n268_ | new_n270_ | new_n267_ | new_n264_ | new_n265_ | new_n224_ | new_n230_ | new_n223_ | new_n219_ | new_n220_ | new_n217_ | new_n218_ | new_n216_ | new_n212_ | new_n213_ | new_n252_ | new_n253_ | new_n247_ | new_n248_ | po41 | new_n240_ | new_n152_ | new_n231_ | new_n150_;
  assign po36 = new_n181_ | new_n192_ | new_n184_ | new_n196_ | new_n199_ | new_n197_ | new_n139_ | new_n153_ | new_n142_ | new_n202_ | new_n141_ | new_n206_ | new_n148_ | new_n310_ | new_n155_ | new_n158_ | new_n311_ | new_n286_ | new_n315_ | new_n297_ | new_n277_ | new_n287_ | new_n289_ | new_n274_ | new_n239_ | new_n240_ | new_n152_ | new_n238_ | new_n229_ | new_n149_ | new_n228_ | new_n208_ | new_n209_ | new_n211_ | po32 | new_n224_ | new_n213_ | new_n220_ | new_n271_ | new_n266_ | new_n268_ | new_n265_ | new_n256_ | new_n205_ | new_n255_ | new_n250_ | new_n253_ | new_n248_ | new_n242_ | new_n166_;
  assign po37 = new_n170_ | new_n169_ | new_n171_ | new_n173_ | new_n172_ | new_n174_ | new_n176_ | new_n175_ | new_n177_ | new_n179_ | new_n178_ | new_n181_ | new_n180_ | new_n182_ | new_n184_ | new_n183_ | new_n185_ | new_n187_ | new_n186_ | new_n188_ | new_n190_ | new_n189_ | new_n192_ | new_n191_ | new_n193_ | new_n195_ | new_n194_ | new_n196_ | new_n198_ | new_n197_ | new_n199_ | new_n201_ | new_n200_ | new_n202_ | new_n204_ | new_n203_ | new_n206_ | new_n136_ | new_n298_ | new_n137_ | new_n141_ | new_n138_ | new_n143_ | new_n140_ | new_n139_ | new_n142_ | new_n144_ | new_n153_ | new_n146_ | new_n145_ | new_n147_ | new_n151_ | new_n148_ | po21 | new_n154_ | new_n156_ | po20 | new_n310_ | new_n155_ | new_n300_ | new_n159_ | new_n158_ | new_n163_ | new_n258_ | new_n165_ | new_n160_ | new_n162_ | new_n161_ | new_n282_ | new_n236_ | new_n285_ | new_n308_ | new_n286_ | new_n311_ | new_n315_ | new_n314_ | new_n313_ | new_n309_ | new_n312_ | new_n303_ | new_n263_ | new_n302_ | new_n307_ | new_n305_ | new_n306_ | new_n304_ | new_n284_ | new_n299_ | new_n281_ | new_n277_ | new_n301_ | new_n297_ | new_n167_ | new_n296_ | new_n294_ | new_n295_ | new_n293_ | new_n292_ | new_n116_ | new_n291_ | new_n289_ | new_n290_ | new_n288_ | new_n245_ | new_n287_ | new_n244_ | new_n243_ | new_n283_ | new_n239_ | new_n280_ | new_n261_ | new_n278_ | new_n227_ | new_n235_ | new_n275_ | new_n276_ | new_n274_ | new_n272_ | new_n273_ | new_n268_ | new_n266_ | new_n267_ | new_n271_ | new_n269_ | new_n270_ | new_n262_ | new_n260_ | new_n168_ | new_n265_ | new_n205_ | new_n264_ | new_n259_ | new_n257_ | new_n135_ | new_n256_ | new_n254_ | new_n255_ | new_n252_ | new_n253_ | new_n251_ | new_n249_ | new_n250_ | new_n166_ | new_n242_ | new_n164_ | new_n248_ | new_n226_ | new_n247_ | new_n152_ | new_n234_ | new_n150_ | new_n233_ | new_n231_ | new_n232_ | new_n238_ | new_n157_ | new_n237_ | new_n241_ | po41 | new_n240_ | new_n229_ | new_n230_ | new_n228_ | new_n225_ | new_n149_ | new_n224_ | new_n221_ | new_n223_ | new_n220_ | new_n218_ | new_n219_ | new_n214_ | new_n212_ | new_n213_ | new_n217_ | new_n215_ | new_n216_ | po32 | new_n209_ | new_n211_ | new_n208_ | new_n207_ | (pi18 & pi19 & pi20 & pi21 & pi26 & pi30);
  assign po38 = (~pi00 & ((((~pi18 & ~pi19 & pi20 & pi21 & ~pi29 & pi30) | (pi18 & pi19 & ~pi20 & ~pi21 & pi29 & ~pi30)) & (pi22 | pi25)) | (~pi21 & (pi20 ? (pi29 ? ((~pi30 & (pi18 ? ((~pi19 & ~pi28 & pi26) | (~pi27 & ~pi04 & pi19 & pi28)) : (pi19 ? (pi22 & (pi28 | (~pi28 & ~pi05))) : (~pi28 & pi23)))) | (pi18 & pi19 & ~pi28 & pi30 & ~pi27 & ~pi05)) : ((pi18 & ((~pi19 & pi28 & pi30 & pi26 & pi11) | (pi19 & pi03 & pi27))) | (~pi18 & ~pi19 & pi28 & pi30 & ~pi03 & pi02))) : (pi18 ? (pi19 & pi26 & (pi28 ? (~pi29 & pi30) : (pi29 & ~pi30))) : (~pi19 & ~pi03 & ((~pi28 & pi29 & ~pi30 & ~pi05) | (pi28 & ~pi29 & pi30 & ~pi02)))))) | (pi21 & ~pi29 & pi30 & ((~pi18 & (pi19 ? (pi28 | (pi20 & pi22 & ~pi28 & ~pi05 & ~pi15)) : (pi20 & pi26))) | (~pi28 & ~pi05 & ~pi15 & pi18 & ~pi19 & pi20))))) | (~pi01 & ~pi18 & pi19 & ~pi20 & (pi22 | pi23) & ((~pi21 & pi29 & ~pi30) | (~pi29 & pi30 & pi21 & ~pi28))) | new_n222_ | new_n246_ | new_n279_;
  assign po39 = new_n195_ | new_n136_ | new_n200_ | new_n147_ | new_n144_ | po20 | po21 | new_n236_ | new_n302_ | new_n313_ | new_n292_ | new_n167_ | new_n305_ | new_n307_ | new_n213_ | new_n220_ | new_n224_ | new_n230_ | new_n240_ | new_n231_ | new_n152_ | new_n239_ | new_n271_ | new_n274_ | new_n265_ | new_n268_ | new_n248_ | new_n253_;
  assign po40 = new_n237_ | new_n257_ | new_n135_ | new_n244_ | new_n204_ | new_n245_ | new_n313_;
  assign po41 = pi30 & ~pi29 & ~pi28 & pi22 & pi21 & pi20 & pi19 & ~pi18 & ~pi15 & pi00 & ~pi05;
  assign po43 = new_n116_ | new_n293_;
  assign new_n135_ = pi30 & ~pi29 & ~pi28 & pi25 & pi21 & pi20 & ~pi19 & pi18 & pi05 & pi10;
  assign new_n136_ = ~pi30 & pi29 & pi28 & pi26 & ~pi21 & ~pi20 & pi18 & pi19;
  assign new_n137_ = pi30 & ~pi29 & pi28 & pi26 & ~pi21 & ~pi20 & pi19 & pi18 & pi00 & ~pi11;
  assign new_n138_ = pi30 & ~pi29 & pi28 & pi26 & ~pi21 & ~pi20 & pi19 & pi18 & pi00 & pi11;
  assign new_n139_ = ~pi30 & pi29 & ~pi28 & pi26 & ~pi21 & ~pi20 & pi19 & pi00 & pi18;
  assign new_n140_ = pi30 & ~pi29 & ~pi28 & pi26 & ~pi21 & ~pi20 & pi18 & pi19;
  assign new_n141_ = ~pi30 & ~pi29 & pi28 & pi26 & ~pi21 & ~pi20 & pi18 & pi19;
  assign new_n142_ = ~pi30 & pi29 & pi25 & ~pi21 & ~pi20 & pi19 & pi18 & ~pi11 & pi00 & pi10;
  assign new_n143_ = pi30 & pi29 & ~pi28 & pi26 & ~pi21 & ~pi20 & pi18 & pi19;
  assign new_n144_ = pi30 & pi29 & pi25 & ~pi21 & ~pi20 & pi18 & pi19;
  assign new_n145_ = pi30 & ~pi29 & pi25 & ~pi21 & ~pi20 & pi19 & pi10 & pi18;
  assign new_n146_ = pi30 & ~pi29 & pi25 & ~pi21 & ~pi20 & pi19 & ~pi10 & pi18;
  assign new_n147_ = pi30 & pi29 & pi22 & ~pi21 & ~pi20 & pi18 & pi19;
  assign new_n148_ = ~pi30 & pi29 & pi22 & ~pi21 & ~pi20 & pi19 & pi00 & pi18;
  assign new_n149_ = pi30 & ~pi29 & ~pi28 & pi24 & pi21 & ~pi18 & pi19;
  assign new_n150_ = pi30 & ~pi29 & pi28 & pi21 & pi19 & pi00 & ~pi18;
  assign new_n151_ = pi30 & ~pi29 & pi22 & ~pi21 & ~pi20 & pi18 & pi19;
  assign new_n152_ = ~pi30 & pi29 & pi28 & pi21 & ~pi18 & pi19;
  assign new_n153_ = ~pi30 & pi29 & pi25 & ~pi21 & ~pi20 & pi19 & pi18 & pi11 & pi00 & pi10;
  assign new_n154_ = pi30 & ~pi29 & pi28 & pi26 & ~pi21 & pi20 & ~pi19 & pi18 & pi00 & ~pi11;
  assign new_n155_ = ~pi30 & ~pi29 & pi28 & pi26 & ~pi21 & pi20 & ~pi19 & pi17 & pi18;
  assign new_n156_ = pi30 & ~pi29 & pi28 & pi26 & ~pi21 & pi20 & ~pi19 & pi18 & pi00 & pi11;
  assign new_n157_ = pi30 & pi29 & pi28 & pi21 & ~pi18 & pi19;
  assign new_n158_ = ~pi30 & pi29 & ~pi28 & pi26 & ~pi21 & pi20 & ~pi19 & pi18 & pi00 & pi17;
  assign new_n159_ = pi30 & ~pi29 & ~pi28 & pi26 & ~pi21 & pi20 & ~pi19 & ~pi17 & pi18;
  assign new_n160_ = pi30 & ~pi29 & ~pi28 & pi26 & ~pi21 & pi20 & ~pi19 & pi17 & pi18;
  assign new_n161_ = pi30 & pi23 & ~pi21 & pi20 & pi18 & ~pi19;
  assign new_n162_ = pi30 & pi22 & ~pi21 & pi20 & pi18 & ~pi19;
  assign new_n163_ = pi30 & pi25 & ~pi21 & ~pi20 & ~pi19 & ~pi10 & pi18;
  assign new_n164_ = ~pi30 & ~pi29 & pi28 & pi22 & pi21 & pi20 & pi19 & ~pi18 & pi08 & pi16;
  assign new_n165_ = pi30 & pi25 & ~pi21 & ~pi20 & ~pi19 & pi10 & pi18;
  assign new_n166_ = ~pi30 & ~pi29 & pi28 & pi22 & pi21 & pi20 & pi19 & ~pi18 & ~pi07 & ~pi16;
  assign new_n167_ = pi30 & pi29 & ~pi28 & ~pi21 & pi20 & ~pi18 & ~pi19;
  assign new_n168_ = pi28 & pi21 & pi20 & ~pi19 & pi18 & pi08 & pi16;
  assign new_n169_ = ~pi37 & ~pi36 & ~pi35 & ~pi34 & ~pi33 & ~pi32 & ~pi31 & ~pi30 & pi29 & pi23 & pi21 & ~pi20 & ~pi18 & ~pi19;
  assign new_n170_ = pi37 & ~pi36 & ~pi35 & ~pi34 & ~pi33 & ~pi32 & ~pi31 & ~pi30 & pi29 & pi23 & pi21 & ~pi20 & ~pi18 & ~pi19;
  assign new_n171_ = pi36 & ~pi35 & ~pi34 & ~pi33 & ~pi32 & ~pi31 & ~pi30 & pi29 & pi23 & pi21 & ~pi20 & ~pi18 & ~pi19;
  assign new_n172_ = pi35 & ~pi34 & ~pi33 & ~pi32 & ~pi31 & ~pi30 & pi29 & pi23 & pi21 & ~pi20 & ~pi18 & ~pi19;
  assign new_n173_ = pi34 & ~pi33 & ~pi32 & ~pi31 & ~pi30 & pi29 & pi23 & pi21 & ~pi20 & ~pi18 & ~pi19;
  assign new_n174_ = pi33 & ~pi32 & ~pi31 & ~pi30 & pi29 & pi23 & pi21 & ~pi20 & ~pi18 & ~pi19;
  assign new_n175_ = pi32 & ~pi31 & ~pi30 & pi29 & pi23 & pi21 & ~pi20 & ~pi18 & ~pi19;
  assign new_n176_ = pi31 & ~pi30 & pi29 & pi23 & pi21 & ~pi20 & ~pi18 & ~pi19;
  assign new_n177_ = pi30 & ~pi29 & pi23 & pi21 & ~pi20 & ~pi18 & ~pi19;
  assign new_n178_ = ~pi44 & pi43 & ~pi42 & ~pi41 & ~pi40 & ~pi39 & ~pi38 & ~pi30 & pi29 & ~pi28 & pi22 & pi21 & ~pi20 & ~pi19 & ~pi09 & ~pi18;
  assign new_n179_ = ~pi44 & ~pi43 & ~pi42 & ~pi41 & ~pi40 & ~pi39 & ~pi38 & ~pi30 & pi29 & ~pi28 & pi22 & pi21 & ~pi20 & ~pi19 & ~pi09 & ~pi18;
  assign new_n180_ = pi44 & ~pi43 & ~pi42 & ~pi41 & ~pi40 & ~pi39 & ~pi38 & ~pi30 & pi29 & ~pi28 & pi22 & pi21 & ~pi20 & ~pi19 & ~pi09 & ~pi18;
  assign new_n181_ = ~pi42 & ~pi41 & pi40 & ~pi39 & ~pi38 & ~pi30 & pi29 & ~pi28 & pi22 & pi21 & ~pi20 & ~pi19 & ~pi09 & ~pi18;
  assign new_n182_ = pi30 & pi28 & pi22 & pi21 & ~pi20 & ~pi18 & ~pi19;
  assign new_n183_ = pi30 & pi29 & ~pi28 & pi22 & pi21 & ~pi20 & ~pi18 & ~pi19;
  assign new_n184_ = pi42 & ~pi41 & pi39 & ~pi38 & ~pi30 & pi29 & ~pi28 & pi22 & pi21 & ~pi20 & ~pi19 & ~pi09 & ~pi18;
  assign new_n185_ = ~pi42 & ~pi41 & pi39 & ~pi38 & ~pi30 & pi29 & ~pi28 & pi22 & pi21 & ~pi20 & ~pi19 & ~pi09 & ~pi18;
  assign new_n186_ = pi42 & ~pi41 & ~pi39 & ~pi38 & ~pi30 & pi29 & ~pi28 & pi22 & pi21 & ~pi20 & ~pi19 & ~pi09 & ~pi18;
  assign new_n187_ = pi41 & ~pi38 & ~pi30 & pi29 & ~pi28 & pi22 & pi21 & ~pi20 & ~pi19 & ~pi09 & ~pi18;
  assign new_n188_ = pi38 & ~pi30 & pi29 & ~pi28 & pi22 & pi21 & ~pi20 & ~pi19 & ~pi09 & ~pi18;
  assign new_n189_ = pi39 & ~pi33 & ~pi31 & pi30 & ~pi29 & ~pi28 & pi22 & pi21 & ~pi20 & ~pi19 & pi09 & ~pi18;
  assign new_n190_ = ~pi39 & ~pi33 & ~pi31 & pi30 & ~pi29 & ~pi28 & pi22 & pi21 & ~pi20 & ~pi19 & pi09 & ~pi18;
  assign new_n191_ = pi31 & pi30 & ~pi29 & ~pi28 & pi22 & pi21 & ~pi20 & ~pi19 & pi09 & ~pi18;
  assign new_n192_ = pi33 & pi30 & ~pi29 & ~pi28 & pi22 & pi21 & ~pi20 & ~pi19 & pi09 & ~pi18;
  assign new_n193_ = pi30 & ~pi29 & ~pi28 & pi22 & pi21 & ~pi20 & ~pi19 & ~pi09 & ~pi18;
  assign new_n194_ = ~pi30 & pi29 & ~pi28 & pi27 & ~pi21 & pi20 & pi18 & pi19;
  assign new_n195_ = pi30 & ~pi29 & pi27 & ~pi21 & pi20 & pi18 & pi19;
  assign new_n196_ = ~pi30 & ~pi29 & pi27 & ~pi21 & pi20 & pi19 & pi18 & pi00 & pi03;
  assign new_n197_ = ~pi30 & ~pi29 & pi27 & ~pi21 & pi20 & pi19 & ~pi03 & pi18;
  assign new_n198_ = pi30 & pi29 & pi28 & ~pi27 & ~pi21 & pi20 & pi18 & pi19;
  assign new_n199_ = ~pi30 & pi29 & pi28 & ~pi27 & ~pi21 & pi20 & pi19 & pi18 & ~pi00 & ~pi04;
  assign new_n200_ = ~pi30 & pi29 & pi28 & ~pi27 & ~pi21 & pi20 & pi19 & pi04 & pi18;
  assign new_n201_ = pi30 & ~pi29 & pi28 & ~pi27 & ~pi21 & pi20 & pi18 & pi19;
  assign new_n202_ = ~pi30 & ~pi29 & pi28 & ~pi27 & ~pi21 & pi20 & pi18 & pi19;
  assign new_n203_ = pi30 & pi29 & ~pi28 & ~pi27 & ~pi21 & pi20 & pi19 & pi18 & pi00 & ~pi05;
  assign new_n204_ = pi30 & pi29 & ~pi28 & ~pi27 & ~pi21 & pi20 & pi19 & pi05 & pi18;
  assign new_n205_ = pi28 & pi21 & pi20 & ~pi19 & pi18 & ~pi08 & pi16;
  assign new_n206_ = ~pi30 & pi29 & ~pi28 & ~pi27 & ~pi21 & pi20 & pi18 & pi19;
  assign new_n207_ = ~pi30 & ~pi29 & ~pi28 & pi14 & ~pi27;
  assign new_n208_ = ~pi30 & ~pi29 & ~pi28 & ~pi27 & ~pi23 & ~pi21 & pi20 & ~pi19 & ~pi14 & ~pi18;
  assign new_n209_ = ~pi30 & ~pi29 & ~pi28 & ~pi27 & ~pi21 & ~pi20 & ~pi19 & ~pi14 & pi18;
  assign new_n210_ = ~pi30 & ~pi29 & ~pi28 & ~pi27 & pi21 & pi13 & ~pi14;
  assign new_n211_ = ~pi30 & ~pi29 & ~pi28 & ~pi27 & ~pi21 & pi13 & ~pi14;
  assign new_n212_ = pi30 & ~pi29 & pi22 & pi21 & pi20 & ~pi19 & pi00 & ~pi18;
  assign new_n213_ = ~pi30 & pi29 & ~pi26 & pi21 & pi20 & ~pi18 & ~pi19;
  assign new_n214_ = pi30 & pi29 & ~pi26 & pi21 & pi20 & ~pi18 & ~pi19;
  assign new_n215_ = pi25 & pi21 & pi20 & ~pi19 & ~pi10 & ~pi18;
  assign new_n216_ = pi30 & ~pi29 & pi25 & pi21 & pi20 & ~pi19 & ~pi18 & ~pi11 & pi00 & pi10;
  assign new_n217_ = pi30 & ~pi29 & pi25 & pi21 & pi20 & ~pi19 & ~pi18 & pi11 & pi00 & pi10;
  assign new_n218_ = pi30 & ~pi29 & pi26 & pi21 & pi20 & ~pi19 & ~pi18 & pi00 & ~pi11;
  assign new_n219_ = pi30 & ~pi29 & pi26 & pi21 & pi20 & ~pi19 & ~pi18 & pi00 & pi11;
  assign new_n220_ = ~pi30 & pi29 & pi26 & pi21 & pi20 & ~pi18 & ~pi19;
  assign new_n221_ = pi30 & pi29 & pi26 & pi21 & pi20 & ~pi18 & ~pi19;
  assign new_n222_ = pi30 & ~pi29 & pi24 & pi21 & pi20 & ~pi19 & ~pi00 & ~pi18;
  assign new_n223_ = pi30 & ~pi29 & pi24 & pi21 & pi20 & ~pi19 & pi00 & ~pi18;
  assign new_n224_ = ~pi30 & pi29 & pi24 & pi21 & pi20 & ~pi18 & ~pi19;
  assign new_n225_ = pi30 & pi29 & pi24 & pi21 & pi20 & ~pi18 & ~pi19;
  assign new_n226_ = ~pi30 & ~pi29 & pi28 & pi22 & pi21 & pi20 & pi19 & ~pi18 & pi07 & ~pi16;
  assign new_n227_ = pi30 & pi25 & pi21 & ~pi20 & pi19 & pi10 & pi18;
  assign new_n228_ = pi30 & ~pi29 & ~pi28 & pi25 & pi21 & pi19 & pi10 & ~pi18;
  assign new_n229_ = pi30 & ~pi29 & ~pi28 & pi26 & pi21 & ~pi18 & pi19;
  assign new_n230_ = pi30 & ~pi29 & ~pi28 & pi22 & pi21 & ~pi20 & pi19 & pi01 & ~pi18;
  assign new_n231_ = pi30 & ~pi29 & ~pi28 & pi23 & pi21 & ~pi20 & pi19 & pi01 & ~pi18;
  assign new_n232_ = pi30 & ~pi29 & ~pi28 & pi25 & pi21 & pi19 & ~pi10 & ~pi18;
  assign new_n233_ = ~pi30 & pi29 & ~pi28 & pi22 & pi21 & ~pi20 & ~pi18 & pi19;
  assign new_n234_ = ~pi30 & pi29 & ~pi28 & pi23 & pi21 & ~pi20 & ~pi18 & pi19;
  assign new_n235_ = pi30 & pi26 & pi21 & ~pi20 & pi18 & pi19;
  assign new_n236_ = pi30 & ~pi29 & pi28 & pi22 & ~pi21 & pi20 & pi19 & ~pi18 & pi02 & ~pi03;
  assign new_n237_ = pi30 & ~pi29 & ~pi28 & pi22 & pi21 & pi20 & pi19 & pi05 & ~pi18;
  assign new_n238_ = pi30 & ~pi29 & ~pi28 & pi22 & pi21 & pi20 & pi19 & ~pi18 & ~pi05 & pi15;
  assign new_n239_ = ~pi30 & pi29 & pi21 & pi20 & pi18 & pi19;
  assign new_n240_ = ~pi30 & pi29 & ~pi28 & pi22 & pi21 & pi20 & ~pi18 & pi19;
  assign new_n241_ = pi30 & pi29 & ~pi28 & pi22 & pi21 & pi20 & ~pi18 & pi19;
  assign new_n242_ = ~pi30 & ~pi29 & pi28 & pi22 & pi21 & pi20 & pi19 & ~pi18 & ~pi08 & pi16;
  assign new_n243_ = pi30 & pi29 & pi21 & pi20 & pi18 & pi19;
  assign new_n244_ = ~pi30 & pi29 & ~pi28 & ~pi21 & ~pi20 & ~pi19 & pi03 & ~pi18;
  assign new_n245_ = ~pi30 & pi29 & ~pi28 & ~pi21 & ~pi20 & ~pi19 & ~pi18 & ~pi03 & pi05;
  assign new_n246_ = pi30 & ~pi29 & ~pi28 & pi21 & ~pi20 & ~pi19 & ~pi00 & pi18;
  assign new_n247_ = pi30 & ~pi29 & ~pi28 & pi21 & ~pi20 & ~pi19 & pi00 & pi18;
  assign new_n248_ = ~pi30 & pi29 & ~pi28 & pi21 & ~pi20 & pi18 & ~pi19;
  assign new_n249_ = pi30 & pi29 & ~pi28 & pi21 & ~pi20 & pi18 & ~pi19;
  assign new_n250_ = ~pi30 & ~pi29 & pi28 & pi21 & ~pi20 & pi18 & ~pi19;
  assign new_n251_ = pi30 & ~pi29 & pi28 & pi21 & ~pi20 & pi18 & ~pi19;
  assign new_n252_ = pi30 & ~pi29 & ~pi28 & pi22 & pi21 & pi20 & ~pi19 & pi18 & ~pi15 & pi00 & ~pi05;
  assign new_n253_ = ~pi30 & pi29 & ~pi28 & pi22 & pi21 & pi20 & pi18 & ~pi19;
  assign new_n254_ = pi30 & pi29 & ~pi28 & pi22 & pi21 & pi20 & pi18 & ~pi19;
  assign new_n255_ = pi30 & ~pi29 & ~pi28 & pi21 & pi20 & ~pi19 & pi18 & ~pi05 & pi15;
  assign new_n256_ = pi28 & pi21 & pi20 & ~pi19 & pi18 & ~pi07 & ~pi16;
  assign new_n257_ = pi30 & ~pi29 & ~pi28 & ~pi25 & pi21 & pi20 & ~pi19 & pi05 & pi18;
  assign new_n258_ = pi30 & pi22 & ~pi21 & ~pi20 & pi18 & ~pi19;
  assign new_n259_ = pi30 & ~pi29 & ~pi28 & pi25 & pi21 & pi20 & ~pi19 & pi18 & pi05 & ~pi10;
  assign new_n260_ = pi30 & ~pi29 & ~pi28 & pi25 & pi21 & pi20 & ~pi19 & pi18 & ~pi15 & ~pi10 & pi00 & ~pi05;
  assign new_n261_ = pi30 & ~pi29 & pi21 & pi20 & pi19 & pi00 & pi18;
  assign new_n262_ = pi28 & pi21 & pi20 & ~pi19 & pi18 & pi07 & ~pi16;
  assign new_n263_ = pi30 & ~pi29 & pi23 & ~pi21 & ~pi20 & ~pi18 & pi19;
  assign new_n264_ = pi30 & ~pi29 & ~pi28 & pi25 & pi21 & pi20 & ~pi19 & pi18 & ~pi15 & ~pi11 & pi10 & pi00 & ~pi05;
  assign new_n265_ = ~pi30 & pi29 & ~pi28 & pi25 & pi21 & pi20 & ~pi19 & ~pi11 & pi18;
  assign new_n266_ = pi30 & pi29 & ~pi28 & pi25 & pi21 & pi20 & ~pi19 & ~pi11 & pi18;
  assign new_n267_ = pi30 & ~pi29 & ~pi28 & pi25 & pi21 & pi20 & ~pi19 & pi18 & ~pi15 & pi11 & pi10 & pi00 & ~pi05;
  assign new_n268_ = ~pi30 & pi29 & ~pi28 & pi25 & pi21 & pi20 & ~pi19 & pi11 & pi18;
  assign new_n269_ = pi30 & pi29 & ~pi28 & pi25 & pi21 & pi20 & ~pi19 & pi11 & pi18;
  assign new_n270_ = pi30 & ~pi29 & ~pi28 & pi26 & pi21 & pi20 & ~pi19 & pi18 & ~pi15 & ~pi11 & pi00 & ~pi05;
  assign new_n271_ = ~pi30 & pi29 & ~pi28 & pi26 & pi21 & pi20 & ~pi19 & ~pi11 & pi18;
  assign new_n272_ = pi30 & pi29 & ~pi28 & pi26 & pi21 & pi20 & ~pi19 & ~pi11 & pi18;
  assign new_n273_ = pi30 & ~pi29 & ~pi28 & pi26 & pi21 & pi20 & ~pi19 & pi18 & ~pi15 & pi11 & pi00 & ~pi05;
  assign new_n274_ = ~pi30 & pi29 & ~pi28 & pi26 & pi21 & pi20 & ~pi19 & pi11 & pi18;
  assign new_n275_ = pi30 & pi29 & ~pi28 & pi26 & pi21 & pi20 & ~pi19 & pi11 & pi18;
  assign new_n276_ = pi30 & pi22 & pi21 & ~pi20 & pi18 & pi19;
  assign new_n277_ = ~pi30 & ~pi29 & pi28 & ~pi21 & pi20 & ~pi18 & ~pi19;
  assign new_n278_ = pi30 & pi25 & pi21 & ~pi20 & pi19 & ~pi10 & pi18;
  assign new_n279_ = pi30 & ~pi29 & pi24 & pi21 & pi20 & pi19 & ~pi00 & pi18;
  assign new_n280_ = pi30 & pi22 & pi21 & pi20 & pi18 & pi19;
  assign new_n281_ = pi30 & ~pi29 & pi28 & ~pi21 & pi20 & ~pi19 & ~pi18 & ~pi06 & ~pi02 & ~pi03;
  assign new_n282_ = pi30 & ~pi29 & pi28 & pi22 & ~pi21 & pi20 & pi19 & ~pi18 & ~pi02 & ~pi03;
  assign new_n283_ = pi30 & ~pi29 & ~pi28 & ~pi21 & ~pi20 & ~pi18 & ~pi19;
  assign new_n284_ = pi30 & ~pi29 & pi28 & ~pi21 & pi20 & ~pi19 & ~pi18 & pi03 & pi06;
  assign new_n285_ = pi30 & pi29 & pi28 & pi22 & ~pi21 & pi20 & ~pi18 & pi19;
  assign new_n286_ = ~pi30 & pi29 & pi28 & pi22 & ~pi21 & pi20 & pi19 & pi00 & ~pi18;
  assign new_n287_ = ~pi30 & pi29 & ~pi28 & ~pi21 & ~pi20 & ~pi19 & ~pi18 & ~pi05 & pi00 & ~pi03;
  assign new_n288_ = pi30 & pi29 & ~pi28 & ~pi21 & ~pi20 & ~pi18 & ~pi19;
  assign new_n289_ = ~pi30 & ~pi29 & pi28 & ~pi21 & ~pi20 & ~pi18 & ~pi19;
  assign new_n290_ = pi30 & ~pi29 & pi28 & ~pi21 & ~pi20 & ~pi19 & ~pi18 & ~pi02 & ~pi03;
  assign new_n291_ = pi30 & ~pi29 & pi28 & ~pi21 & ~pi20 & ~pi19 & ~pi18 & ~pi03 & pi00 & pi02;
  assign new_n292_ = ~pi30 & pi29 & pi28 & ~pi21 & ~pi20 & ~pi18 & ~pi19;
  assign new_n293_ = pi30 & ~pi29 & pi24 & ~pi21 & pi20 & ~pi18 & ~pi19;
  assign new_n294_ = ~pi30 & pi29 & pi24 & ~pi21 & pi20 & ~pi18 & ~pi19;
  assign new_n295_ = pi30 & ~pi29 & pi26 & ~pi21 & pi20 & ~pi18 & ~pi19;
  assign new_n296_ = pi30 & ~pi29 & ~pi28 & pi23 & ~pi21 & pi20 & ~pi18 & ~pi19;
  assign new_n297_ = ~pi30 & pi29 & ~pi28 & pi23 & ~pi21 & pi20 & ~pi19 & pi00 & ~pi18;
  assign new_n298_ = pi30 & ~pi29 & ~pi28 & ~pi27 & ~pi21 & pi20 & pi18 & pi19;
  assign new_n299_ = pi30 & ~pi29 & pi28 & ~pi21 & pi20 & ~pi19 & ~pi18 & pi06 & ~pi02 & ~pi03;
  assign new_n300_ = ~pi30 & pi29 & ~pi28 & pi26 & ~pi21 & pi20 & ~pi19 & pi17 & pi18;
  assign new_n301_ = pi30 & ~pi29 & pi28 & ~pi21 & pi20 & ~pi19 & ~pi18 & pi03 & ~pi06;
  assign new_n302_ = ~pi30 & pi29 & pi23 & ~pi21 & ~pi20 & pi19 & pi01 & ~pi18;
  assign new_n303_ = pi30 & ~pi29 & ~pi28 & pi22 & ~pi21 & pi20 & ~pi18 & pi19;
  assign new_n304_ = pi30 & ~pi29 & pi28 & ~pi21 & pi20 & ~pi19 & ~pi18 & ~pi03 & pi00 & ~pi02;
  assign new_n305_ = ~pi30 & pi29 & pi28 & ~pi21 & pi20 & ~pi18 & ~pi19;
  assign new_n306_ = pi30 & ~pi29 & pi22 & ~pi21 & ~pi20 & ~pi18 & pi19;
  assign new_n307_ = ~pi30 & pi29 & pi22 & ~pi21 & ~pi20 & pi19 & pi01 & ~pi18;
  assign new_n308_ = pi30 & ~pi29 & pi28 & pi22 & ~pi21 & pi20 & pi19 & pi03 & ~pi18;
  assign new_n309_ = pi30 & ~pi29 & ~pi28 & pi23 & ~pi21 & pi20 & ~pi18 & pi19;
  assign new_n310_ = ~pi30 & pi29 & ~pi28 & pi26 & ~pi21 & pi20 & ~pi19 & pi18 & pi00 & ~pi17;
  assign new_n311_ = ~pi30 & ~pi29 & pi28 & pi22 & ~pi21 & pi20 & ~pi18 & pi19;
  assign new_n312_ = pi30 & ~pi29 & ~pi28 & pi26 & ~pi21 & pi20 & ~pi18 & pi19;
  assign new_n313_ = ~pi30 & pi29 & ~pi28 & pi22 & ~pi21 & pi20 & pi19 & pi05 & ~pi18;
  assign new_n314_ = pi30 & pi29 & ~pi28 & pi22 & ~pi21 & pi20 & ~pi18 & pi19;
  assign new_n315_ = ~pi30 & pi29 & ~pi28 & pi22 & ~pi21 & pi20 & pi19 & ~pi18 & pi00 & ~pi05;
  assign po24 = new_n116_;
  assign po44 = new_n116_;
  assign po02 = 1'b0;
  assign po42 = 1'b0;
endmodule


