// Benchmark "apex6" written by ABC on Thu Mar 19 13:02:36 2020

module apex6 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47,
    po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71,
    po72, po73, po74, po75, po76, po77, po78, po79, po80, po81, po82, po83,
    po84, po85, po86, po87, po88, po89, po90, po91, po92, po93, po94, po95,
    po96, po97, po98  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46,
    po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58,
    po59, po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70,
    po71, po72, po73, po74, po75, po76, po77, po78, po79, po80, po81, po82,
    po83, po84, po85, po86, po87, po88, po89, po90, po91, po92, po93, po94,
    po95, po96, po97, po98;
  wire new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_;
  assign po00 = ~pi072 | pi075;
  assign po01 = pi073 | (~pi001 & new_n334_ & new_n335_);
  assign po02 = new_n336_ & ~pi073;
  assign po03 = (pi081 & po45) | (~pi038 & pi077);
  assign po04 = (pi040 & new_n337_) | (pi008 & new_n338_);
  assign po05 = (pi041 & new_n337_) | (pi009 & new_n338_);
  assign po06 = (pi042 & new_n337_) | (pi010 & new_n338_);
  assign po07 = (pi043 & new_n337_) | (pi011 & new_n338_);
  assign po08 = (pi044 & new_n337_) | (pi012 & new_n338_);
  assign po09 = (pi045 & new_n337_) | (pi013 & new_n338_);
  assign po10 = (pi046 & new_n337_) | (pi014 & new_n338_);
  assign po11 = (pi047 & new_n337_) | (pi015 & new_n338_);
  assign po12 = (pi048 & new_n339_) | (pi008 & new_n340_);
  assign po13 = (pi049 & new_n339_) | (pi009 & new_n340_);
  assign po14 = (pi050 & new_n339_) | (pi010 & new_n340_);
  assign po15 = (pi051 & new_n339_) | (pi011 & new_n340_);
  assign po16 = (pi052 & new_n339_) | (pi012 & new_n340_);
  assign po17 = (pi053 & new_n339_) | (pi013 & new_n340_);
  assign po18 = (pi054 & new_n339_) | (pi014 & new_n340_);
  assign po19 = (pi055 & new_n339_) | (pi015 & new_n340_);
  assign po20 = (pi056 & new_n341_) | (pi018 & new_n342_);
  assign po21 = (pi057 & new_n341_) | (pi019 & new_n342_);
  assign po22 = (pi058 & new_n341_) | (pi020 & new_n342_);
  assign po23 = (pi059 & new_n341_) | (pi021 & new_n342_);
  assign po24 = (pi060 & new_n341_) | (pi022 & new_n342_);
  assign po25 = (pi061 & new_n341_) | (pi023 & new_n342_);
  assign po26 = (pi062 & new_n341_) | (pi024 & new_n342_);
  assign po27 = (pi063 & new_n341_) | (pi025 & new_n342_);
  assign po28 = (pi064 & new_n343_) | (pi018 & new_n344_);
  assign po29 = (pi065 & new_n343_) | (pi019 & new_n344_);
  assign po30 = (pi066 & new_n343_) | (pi020 & new_n344_);
  assign po31 = (pi067 & new_n343_) | (pi021 & new_n344_);
  assign po32 = (pi068 & new_n343_) | (pi022 & new_n344_);
  assign po33 = (pi069 & new_n343_) | (pi023 & new_n344_);
  assign po34 = (pi070 & new_n343_) | (pi024 & new_n344_);
  assign po35 = (pi071 & new_n343_) | (pi025 & new_n344_);
  assign po36 = pi073 | new_n345_;
  assign po37 = pi038 | (pi083 & new_n346_);
  assign po38 = new_n347_ & ~pi073;
  assign po39 = new_n348_ & ~pi073;
  assign po40 = pi076 ? new_n349_ : (~new_n350_ & new_n351_);
  assign po41 = (pi077 & new_n352_) | (pi076 & ~pi077 & new_n351_ & ~new_n350_);
  assign po42 = new_n354_ & pi000 & new_n353_;
  assign po43 = (~pi079 & new_n355_) | (~pi075 & pi079 & new_n356_);
  assign po44 = (pi080 & new_n357_) | (pi079 & ~pi080 & new_n355_);
  assign po45 = ~pi038 & pi082;
  assign po46 = pi036 & ~pi038;
  assign po47 = new_n358_ & ~pi073;
  assign po48 = new_n359_ & ~pi073;
  assign po49 = new_n360_ & ~pi073;
  assign po50 = (~pi073 & pi086 & new_n345_) | (~pi086 & ~po36);
  assign po51 = (pi087 & new_n361_ & ~pi073) | (pi086 & ~pi087 & ~po36);
  assign po52 = pi088 ? (new_n362_ & ~pi073) : new_n363_;
  assign po53 = (pi088 & ~pi089 & new_n363_) | (pi089 & new_n364_ & ~pi073);
  assign po54 = (new_n365_ & pi090 & ~pi073) | (pi088 & pi089 & ~pi090 & new_n363_);
  assign po55 = new_n366_ & ~pi073;
  assign po56 = new_n367_ & ~pi073;
  assign po57 = (pi094 & new_n369_) | (pi093 & new_n368_);
  assign po58 = (pi095 & new_n369_) | (pi094 & new_n368_);
  assign po59 = (pi096 & new_n369_) | (pi095 & new_n368_);
  assign po60 = (pi097 & new_n369_) | (pi096 & new_n368_);
  assign po61 = (pi098 & new_n369_) | (pi097 & new_n368_);
  assign po62 = (pi099 & new_n369_) | (pi098 & new_n368_);
  assign po63 = (pi100 & new_n369_) | (pi099 & new_n368_);
  assign po64 = (pi100 & new_n368_) | (pi005 & new_n369_);
  assign po65 = (pi102 & new_n371_) | (pi101 & new_n370_);
  assign po66 = (pi103 & new_n371_) | (pi102 & new_n370_);
  assign po67 = (pi104 & new_n371_) | (pi103 & new_n370_);
  assign po68 = (pi105 & new_n371_) | (pi104 & new_n370_);
  assign po69 = (pi106 & new_n371_) | (pi105 & new_n370_);
  assign po70 = (pi107 & new_n371_) | (pi106 & new_n370_);
  assign po71 = (pi108 & new_n371_) | (pi107 & new_n370_);
  assign po72 = (pi108 & new_n370_) | (pi005 & new_n371_);
  assign po73 = new_n372_ & ~pi073;
  assign po74 = (new_n374_ & pi057) | (new_n373_ & new_n375_);
  assign po75 = (new_n374_ & pi058) | (new_n373_ & new_n376_);
  assign po76 = (new_n378_ & new_n379_) | (new_n374_ & pi059) | (new_n377_ & pi043);
  assign po77 = (new_n380_ & new_n379_) | (new_n374_ & pi060) | (new_n377_ & pi044);
  assign po78 = (new_n381_ & new_n379_) | (new_n374_ & pi061) | (new_n377_ & pi045);
  assign po79 = (new_n382_ & new_n379_) | (new_n374_ & pi062) | (new_n377_ & pi046);
  assign po80 = new_n383_ & ~pi073;
  assign po81 = (new_n384_ & new_n379_) | (new_n374_ & pi064) | (new_n377_ & pi048);
  assign po82 = (new_n374_ & pi065) | (new_n373_ & new_n385_);
  assign po83 = ~pi073 & new_n386_;
  assign po84 = new_n387_ & ~pi073;
  assign po85 = new_n388_ & ~pi073;
  assign po86 = (new_n389_ & new_n379_) | (new_n377_ & pi053) | (new_n374_ & pi069);
  assign po87 = (new_n374_ & pi070) | (new_n377_ & pi054) | (new_n390_ & new_n379_);
  assign po88 = (new_n374_ & pi071) | (new_n373_ & new_n391_);
  assign po89 = ~pi125 & new_n392_;
  assign po90 = pi126 ? po89 : new_n351_;
  assign po91 = (pi127 & new_n393_) | (pi126 & ~pi127 & new_n351_);
  assign po92 = pi128 ? new_n395_ : (new_n351_ & new_n394_);
  assign po93 = pi129 ? new_n397_ : (new_n396_ & new_n392_);
  assign po94 = (pi130 & new_n398_) | (new_n351_ & ~new_n399_);
  assign po95 = pi131 ? new_n400_ : (~new_n399_ & new_n351_);
  assign po96 = (new_n402_ & pi132) | (new_n401_ & ~pi132 & new_n392_);
  assign po97 = (pi133 & new_n403_) | (new_n401_ & pi132 & ~pi133 & new_n392_);
  assign po98 = new_n354_ & pi000 & new_n404_;
  assign new_n334_ = ~pi002 & ~pi003;
  assign new_n335_ = pi039 | (pi083 & new_n346_);
  assign new_n336_ = (pi075 & pi037 & new_n408_) | (~pi075 & new_n406_ & ~pi072) | (new_n405_ & ~pi089 & ~pi090 & new_n407_);
  assign new_n337_ = new_n409_ & ~pi073;
  assign new_n338_ = ~pi073 & ~new_n409_;
  assign new_n339_ = new_n410_ & ~pi073;
  assign new_n340_ = ~pi073 & ~new_n410_;
  assign new_n341_ = new_n411_ & ~pi073;
  assign new_n342_ = ~pi073 & ~new_n411_;
  assign new_n343_ = new_n412_ & ~pi073;
  assign new_n344_ = ~pi073 & ~new_n412_;
  assign new_n345_ = new_n334_ & pi072 & ~pi001;
  assign new_n346_ = pi092 & ~pi072 & pi091;
  assign new_n347_ = (new_n415_ & pi074) | (new_n414_ & pi083) | (new_n413_ & new_n416_ & ~pi072 & ~pi074);
  assign new_n348_ = new_n419_ | (pi075 & new_n417_) | (~pi032 & ~pi033 & ~new_n418_);
  assign new_n349_ = po89 | (new_n350_ & new_n392_);
  assign new_n350_ = pi133 | new_n420_ | pi132 | ~pi130 | pi131;
  assign new_n351_ = pi125 & new_n392_;
  assign new_n352_ = new_n349_ | (~pi076 & new_n392_);
  assign new_n353_ = po46 | (~pi038 & pi078);
  assign new_n354_ = ~pi081 | ~pi082;
  assign new_n355_ = (new_n421_ & ~pi038) | (po46 & pi078 & ~pi032 & ~pi033 & ~pi034 & ~pi035);
  assign new_n356_ = po89 | (~pi038 & new_n422_);
  assign new_n357_ = (~pi079 & ~pi038) | (~pi075 & new_n356_);
  assign new_n358_ = pi083 | (~pi072 & ~new_n423_);
  assign new_n359_ = (pi084 & new_n426_) | (~new_n424_ & ~new_n425_ & ~pi084 & ~pi089 & ~pi090 & ~pi072);
  assign new_n360_ = pi085 ^ ~new_n427_;
  assign new_n361_ = ~pi086 | new_n345_;
  assign new_n362_ = ~pi087 | new_n361_;
  assign new_n363_ = ~po36 & pi087 & pi086;
  assign new_n364_ = ~pi088 | new_n362_;
  assign new_n365_ = ~pi089 | new_n364_;
  assign new_n366_ = pi091 ^ ~new_n428_;
  assign new_n367_ = (pi092 & new_n429_) | (~new_n428_ & pi091 & ~pi092);
  assign new_n368_ = new_n430_ & ~pi073;
  assign new_n369_ = ~pi073 & ~new_n430_;
  assign new_n370_ = new_n431_ & ~pi073;
  assign new_n371_ = ~pi073 & ~new_n431_;
  assign new_n372_ = (new_n432_ & pi040) | (pi003 & pi056) | (new_n334_ & new_n433_);
  assign new_n373_ = ~pi003 & ~pi073;
  assign new_n374_ = pi003 & ~pi073;
  assign new_n375_ = (pi094 & new_n436_) | (pi111 & new_n435_) | (pi002 & pi041) | (pi110 & new_n434_);
  assign new_n376_ = (pi095 & new_n436_) | (pi112 & new_n435_) | (pi002 & pi042) | (pi111 & new_n434_);
  assign new_n377_ = pi002 & new_n373_;
  assign new_n378_ = (pi113 & new_n438_) | (pi001 & pi096) | (pi112 & new_n437_);
  assign new_n379_ = ~pi002 & new_n373_;
  assign new_n380_ = (pi114 & new_n438_) | (pi001 & pi097) | (pi113 & new_n437_);
  assign new_n381_ = (pi115 & new_n438_) | (pi001 & pi098) | (pi114 & new_n437_);
  assign new_n382_ = (pi116 & new_n438_) | (pi001 & pi099) | (pi115 & new_n437_);
  assign new_n383_ = (new_n432_ & pi047) | (new_n334_ & new_n439_) | (pi003 & pi063);
  assign new_n384_ = (pi118 & new_n438_) | (pi001 & pi101) | (pi117 & new_n437_);
  assign new_n385_ = (pi102 & new_n436_) | (pi119 & new_n435_) | (pi002 & pi049) | (pi118 & new_n434_);
  assign new_n386_ = (pi003 & pi066) | (pi050 & new_n432_) | (new_n440_ & new_n334_);
  assign new_n387_ = (pi003 & pi067) | (pi051 & new_n432_) | (new_n334_ & new_n441_);
  assign new_n388_ = (pi003 & pi068) | (pi052 & new_n432_) | (new_n334_ & new_n442_);
  assign new_n389_ = (pi123 & new_n438_) | (pi001 & pi106) | (pi122 & new_n437_);
  assign new_n390_ = (pi124 & new_n438_) | (pi001 & pi107) | (pi123 & new_n437_);
  assign new_n391_ = (pi108 & new_n436_) | (pi002 & pi055) | (pi124 & new_n434_);
  assign new_n392_ = ~pi036 & ~pi038;
  assign new_n393_ = po89 | (~pi126 & new_n392_);
  assign new_n394_ = pi126 & pi127;
  assign new_n395_ = new_n393_ | (~pi127 & new_n392_);
  assign new_n396_ = new_n394_ & pi125 & pi128;
  assign new_n397_ = new_n393_ | (new_n443_ & new_n392_);
  assign new_n398_ = po89 | (new_n420_ & new_n392_);
  assign new_n399_ = pi130 | new_n420_;
  assign new_n400_ = po89 | (new_n399_ & new_n392_);
  assign new_n401_ = ~new_n399_ & pi125 & pi131;
  assign new_n402_ = new_n400_ | (~pi131 & new_n392_);
  assign new_n403_ = new_n400_ | (new_n392_ & new_n444_);
  assign new_n404_ = (pi078 & po46) | (~pi038 & pi134);
  assign new_n405_ = pi087 ? (~pi088 & new_n445_) : (pi088 & new_n446_);
  assign new_n406_ = (new_n447_ & pi083) | (new_n448_ & pi109 & new_n416_);
  assign new_n407_ = ~po00 | (~pi075 & ~new_n448_ & new_n416_);
  assign new_n408_ = pi028 ? (~pi079 & pi080) : (pi079 & ~pi080);
  assign new_n409_ = ~pi007 | pi016;
  assign new_n410_ = ~pi007 | ~pi016;
  assign new_n411_ = ~pi017 | pi026;
  assign new_n412_ = ~pi017 | ~pi026;
  assign new_n413_ = (new_n448_ & pi109) | (~pi090 & new_n405_ & ~new_n448_ & ~pi089);
  assign new_n414_ = new_n346_ | (new_n450_ & pi074) | (new_n449_ & ~pi072 & ~pi074);
  assign new_n415_ = pi072 | (~new_n413_ & new_n416_);
  assign new_n416_ = ~pi083 | (~pi091 & ~pi092);
  assign new_n417_ = ~pi079 | ~pi080;
  assign new_n418_ = ~pi036 | ~pi078 | pi034 | pi035;
  assign new_n419_ = new_n453_ & new_n452_ & new_n451_ & new_n396_ & pi129 & pi134;
  assign new_n420_ = ~new_n394_ | ~pi128 | ~pi129;
  assign new_n421_ = pi075 | new_n419_;
  assign new_n422_ = (~pi078 & new_n460_) | (pi032 & new_n459_) | (new_n418_ & new_n458_) | (new_n457_ & ~pi036) | (new_n454_ & pi035) | (new_n455_ & pi034) | (pi033 & new_n456_);
  assign new_n423_ = new_n425_ | ~new_n461_;
  assign new_n424_ = ~pi031 | (~pi029 & ~pi030);
  assign new_n425_ = ~pi088 | ~pi086 | pi087;
  assign new_n426_ = new_n425_ | pi090 | pi072 | (new_n424_ & ~pi089);
  assign new_n427_ = pi089 | pi072 | new_n425_ | (~pi090 & new_n462_);
  assign new_n428_ = pi072 | (~pi083 & new_n423_);
  assign new_n429_ = new_n428_ | ~pi091;
  assign new_n430_ = ~pi004 | pi006;
  assign new_n431_ = ~pi004 | ~pi006;
  assign new_n432_ = pi002 & ~pi003;
  assign new_n433_ = (pi110 & new_n438_) | (pi001 & pi093) | (pi109 & new_n437_);
  assign new_n434_ = ~pi002 & new_n437_;
  assign new_n435_ = ~pi002 & new_n438_;
  assign new_n436_ = pi001 & ~pi002;
  assign new_n437_ = ~pi001 & new_n463_;
  assign new_n438_ = ~pi001 & ~new_n463_;
  assign new_n439_ = (pi117 & new_n438_) | (pi001 & pi100) | (pi116 & new_n437_);
  assign new_n440_ = (pi120 & new_n438_) | (pi001 & pi103) | (pi119 & new_n437_);
  assign new_n441_ = (pi121 & new_n438_) | (pi001 & pi104) | (pi120 & new_n437_);
  assign new_n442_ = (pi122 & new_n438_) | (pi001 & pi105) | (pi121 & new_n437_);
  assign new_n443_ = ~pi127 | ~pi128;
  assign new_n444_ = ~pi132 | ~pi131;
  assign new_n445_ = pi086 ? pi034 : pi035;
  assign new_n446_ = pi086 ? pi032 : pi033;
  assign new_n447_ = (new_n464_ & pi092) | (~pi027 & pi091 & ~pi092);
  assign new_n448_ = pi084 | pi085;
  assign new_n449_ = (pi028 & pi092) | (~pi027 & pi091);
  assign new_n450_ = (~pi028 & pi092) | (pi027 & pi091);
  assign new_n451_ = new_n465_ & new_n466_;
  assign new_n452_ = pi131 ^ ~pi033;
  assign new_n453_ = ~pi130 ^ ~pi032;
  assign new_n454_ = ~pi125 | ~pi133 | new_n467_;
  assign new_n455_ = ~pi125 | ~pi132 | new_n468_;
  assign new_n456_ = ~pi131 | ~pi134 | new_n469_ | new_n460_;
  assign new_n457_ = new_n468_ | new_n467_;
  assign new_n458_ = new_n469_ | new_n470_;
  assign new_n459_ = new_n460_ | new_n399_ | new_n470_;
  assign new_n460_ = ~pi125 | new_n457_;
  assign new_n461_ = pi089 ? ~new_n472_ : new_n471_;
  assign new_n462_ = ~pi031 | pi029 | pi030;
  assign new_n463_ = pi072 | ~new_n448_;
  assign new_n464_ = pi091 ? ~pi074 : pi028;
  assign new_n465_ = pi035 ^ ~pi133;
  assign new_n466_ = pi132 ^ ~pi034;
  assign new_n467_ = ~pi034 & pi132;
  assign new_n468_ = ~pi035 & pi133;
  assign new_n469_ = new_n420_ | (~pi032 & ~pi130);
  assign new_n470_ = ~pi134 | (~pi033 & pi131);
  assign new_n471_ = ~pi031 | pi090;
  assign new_n472_ = pi090 | ~pi084;
endmodule


